magic
tech sky130A
magscale 1 2
timestamp 1678766716
<< nwell >>
rect -38 315 682 998
<< nmos >>
rect 197 47 227 223
rect 336 47 366 223
rect 475 47 505 223
<< pmos >>
rect 197 351 227 913
rect 336 351 366 913
rect 475 351 505 913
<< ndiff >>
rect 116 171 197 223
rect 116 137 152 171
rect 186 137 197 171
rect 116 103 197 137
rect 116 69 152 103
rect 186 69 197 103
rect 116 47 197 69
rect 227 47 336 223
rect 366 171 475 223
rect 366 137 404 171
rect 438 137 475 171
rect 366 103 475 137
rect 366 69 404 103
rect 438 69 475 103
rect 366 47 475 69
rect 505 171 586 223
rect 505 137 528 171
rect 562 137 586 171
rect 505 103 586 137
rect 505 69 528 103
rect 562 69 586 103
rect 505 48 586 69
rect 505 47 565 48
<< pdiff >>
rect 116 889 197 913
rect 116 855 140 889
rect 174 855 197 889
rect 116 821 197 855
rect 116 787 140 821
rect 174 787 197 821
rect 116 753 197 787
rect 116 719 140 753
rect 174 719 197 753
rect 116 685 197 719
rect 116 651 140 685
rect 174 651 197 685
rect 116 617 197 651
rect 116 583 140 617
rect 174 583 197 617
rect 116 351 197 583
rect 227 889 336 913
rect 227 855 265 889
rect 299 855 336 889
rect 227 821 336 855
rect 227 787 265 821
rect 299 787 336 821
rect 227 753 336 787
rect 227 719 265 753
rect 299 719 336 753
rect 227 685 336 719
rect 227 651 265 685
rect 299 651 336 685
rect 227 617 336 651
rect 227 583 265 617
rect 299 583 336 617
rect 227 351 336 583
rect 366 889 475 913
rect 366 855 403 889
rect 437 855 475 889
rect 366 821 475 855
rect 366 787 403 821
rect 437 787 475 821
rect 366 753 475 787
rect 366 719 403 753
rect 437 719 475 753
rect 366 685 475 719
rect 366 651 403 685
rect 437 651 475 685
rect 366 617 475 651
rect 366 583 403 617
rect 437 583 475 617
rect 366 351 475 583
rect 505 889 586 913
rect 505 855 528 889
rect 562 855 586 889
rect 505 821 586 855
rect 505 787 528 821
rect 562 787 586 821
rect 505 753 586 787
rect 505 719 528 753
rect 562 719 586 753
rect 505 685 586 719
rect 505 651 528 685
rect 562 651 586 685
rect 505 617 586 651
rect 505 583 528 617
rect 562 583 586 617
rect 505 351 586 583
<< ndiffc >>
rect 152 137 186 171
rect 152 69 186 103
rect 404 137 438 171
rect 404 69 438 103
rect 528 137 562 171
rect 528 69 562 103
<< pdiffc >>
rect 140 855 174 889
rect 140 787 174 821
rect 140 719 174 753
rect 140 651 174 685
rect 140 583 174 617
rect 265 855 299 889
rect 265 787 299 821
rect 265 719 299 753
rect 265 651 299 685
rect 265 583 299 617
rect 403 855 437 889
rect 403 787 437 821
rect 403 719 437 753
rect 403 651 437 685
rect 403 583 437 617
rect 528 855 562 889
rect 528 787 562 821
rect 528 719 562 753
rect 528 651 562 685
rect 528 583 562 617
<< psubdiff >>
rect 36 173 116 223
rect 36 139 58 173
rect 92 139 116 173
rect 36 105 116 139
rect 36 71 58 105
rect 92 71 116 105
rect 36 47 116 71
<< nsubdiff >>
rect 36 889 116 913
rect 36 855 58 889
rect 92 855 116 889
rect 36 821 116 855
rect 36 787 58 821
rect 92 787 116 821
rect 36 753 116 787
rect 36 719 58 753
rect 92 719 116 753
rect 36 685 116 719
rect 36 651 58 685
rect 92 651 116 685
rect 36 617 116 651
rect 36 583 58 617
rect 92 583 116 617
rect 36 351 116 583
<< psubdiffcont >>
rect 58 139 92 173
rect 58 71 92 105
<< nsubdiffcont >>
rect 58 855 92 889
rect 58 787 92 821
rect 58 719 92 753
rect 58 651 92 685
rect 58 583 92 617
<< poly >>
rect 197 913 227 939
rect 336 913 366 939
rect 475 913 505 939
rect 197 314 227 351
rect 336 314 366 351
rect 475 314 505 351
rect 63 304 227 314
rect 63 270 79 304
rect 113 270 147 304
rect 181 270 227 304
rect 63 260 227 270
rect 269 304 405 314
rect 269 270 287 304
rect 321 270 355 304
rect 389 270 405 304
rect 269 260 405 270
rect 475 304 609 314
rect 475 270 491 304
rect 525 270 559 304
rect 593 270 609 304
rect 475 260 609 270
rect 197 223 227 260
rect 336 223 366 260
rect 475 223 505 260
rect 197 21 227 47
rect 336 21 366 47
rect 475 21 505 47
<< polycont >>
rect 79 270 113 304
rect 147 270 181 304
rect 287 270 321 304
rect 355 270 389 304
rect 491 270 525 304
rect 559 270 593 304
<< locali >>
rect 0 943 29 977
rect 63 943 121 977
rect 155 943 213 977
rect 247 943 305 977
rect 339 943 397 977
rect 431 943 489 977
rect 523 943 581 977
rect 615 943 644 977
rect 58 889 92 943
rect 58 821 92 855
rect 58 753 92 787
rect 58 685 92 719
rect 58 617 92 651
rect 58 567 92 583
rect 140 889 174 909
rect 140 821 174 855
rect 140 753 174 787
rect 140 685 174 719
rect 140 617 174 651
rect 140 539 174 583
rect 249 889 315 943
rect 249 855 265 889
rect 299 855 315 889
rect 249 821 315 855
rect 249 787 265 821
rect 299 787 315 821
rect 249 753 315 787
rect 249 719 265 753
rect 299 719 315 753
rect 249 685 315 719
rect 249 651 265 685
rect 299 651 315 685
rect 249 617 315 651
rect 249 583 265 617
rect 299 583 315 617
rect 249 582 315 583
rect 403 889 437 909
rect 403 821 437 855
rect 403 753 437 787
rect 403 685 437 719
rect 403 617 437 651
rect 403 539 437 583
rect 140 505 437 539
rect 528 889 562 909
rect 528 821 562 855
rect 528 753 562 787
rect 528 685 562 719
rect 528 617 562 651
rect 528 471 562 583
rect 423 437 562 471
rect 79 304 181 403
rect 113 270 147 304
rect 79 254 181 270
rect 287 304 389 403
rect 321 270 355 304
rect 287 254 389 270
rect 423 212 457 437
rect 491 304 593 403
rect 525 270 559 304
rect 491 254 593 270
rect 58 173 186 190
rect 92 171 186 173
rect 92 139 152 171
rect 58 137 152 139
rect 58 105 186 137
rect 92 103 186 105
rect 92 71 152 103
rect 58 69 152 71
rect 58 17 186 69
rect 404 178 457 212
rect 404 171 438 178
rect 404 103 438 137
rect 404 51 438 69
rect 498 137 528 171
rect 562 137 584 171
rect 498 103 584 137
rect 498 69 528 103
rect 562 69 584 103
rect 498 17 584 69
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 943 63 977
rect 121 943 155 977
rect 213 943 247 977
rect 305 943 339 977
rect 397 943 431 977
rect 489 943 523 977
rect 581 943 615 977
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 977 644 1000
rect 0 943 29 977
rect 63 943 121 977
rect 155 943 213 977
rect 247 943 305 977
rect 339 943 397 977
rect 431 943 489 977
rect 523 943 581 977
rect 615 943 644 977
rect 0 920 644 943
rect 0 17 644 40
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -40 644 -17
<< labels >>
flabel locali s 121 343 155 377 0 FreeSans 240 0 0 0 A1
port 0 nsew signal input
flabel locali s 305 343 339 377 0 FreeSans 240 0 0 0 A2
port 1 nsew signal input
flabel locali s 531 343 565 377 0 FreeSans 240 0 0 0 B1
port 2 nsew signal input
flabel metal1 s 305 -17 339 17 0 FreeSans 240 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 305 943 339 977 0 FreeSans 240 0 0 0 VPWR
port 4 nsew power bidirectional
flabel locali s 528 743 562 777 0 FreeSans 240 0 0 0 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 960
string LEFclass CORE
string LEForigin 0 0
<< end >>
