* NGSPICE file created from thesis_nor2.ext - technology: sky130A

.subckt thesis_nor2 A1 B1 Y VPWR VGND
X0 VGND.t1 B1.t0 Y.t1 VGND sky130_fd_pr__nfet_01v8 ad=0.3608 pd=2.58 as=0.1804 ps=1.29 w=0.88 l=0.15
X1 Y.t0 A1.t0 VGND.t0 VGND sky130_fd_pr__nfet_01v8 ad=0.1804 pd=1.29 as=0.3608 ps=2.58 w=0.88 l=0.15
X2 Y.t2 B1.t1 a_230_351# VPWR.t2 sky130_fd_pr__pfet_01v8 ad=1.1521 pd=6.44 as=0.57605 ps=3.22 w=2.81 l=0.15
X3 a_230_351# A1.t1 VPWR.t1 VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.57605 pd=3.22 as=1.2645 ps=6.52 w=2.81 l=0.15
R0 B1.n0 B1.t1 510.919
R1 B1.n0 B1.t0 200.832
R2 B1 B1.n0 52.922
R3 Y Y.t2 171.524
R4 Y Y.n0 119.12
R5 Y.n0 Y.t1 27.954
R6 Y.n0 Y.t0 27.954
R7 VGND.n0 VGND.t1 117.636
R8 VGND.n0 VGND.t0 88.723
R9 VGND VGND.n0 0.017
R10 A1.n0 A1.t1 510.919
R11 A1.n0 A1.t0 200.832
R12 A1 A1.n0 70.693
R13 VPWR.n23 VPWR.n0 292.5
R14 VPWR.n20 VPWR.t0 203.074
R15 VPWR.t0 VPWR.t2 155.783
R16 VPWR.n22 VPWR.n21 127.045
R17 VPWR.n3 VPWR.n2 92.731
R18 VPWR.n4 VPWR.n1 92.5
R19 VPWR.n15 VPWR.n14 92.5
R20 VPWR.n11 VPWR.n10 92.5
R21 VPWR.n8 VPWR.n7 92.5
R22 VPWR.n18 VPWR.n17 92.5
R23 VPWR.n14 VPWR.n13 34.545
R24 VPWR.n7 VPWR.n6 34.545
R25 VPWR.n21 VPWR.n20 28.978
R26 VPWR.n0 VPWR.t1 12.619
R27 VPWR.n24 VPWR.n23 6.554
R28 VPWR.n22 VPWR.n19 5.012
R29 VPWR.n18 VPWR.n16 5.012
R30 VPWR.n15 VPWR.n12 5.012
R31 VPWR.n11 VPWR.n9 5.012
R32 VPWR.n8 VPWR.n5 5.012
R33 VPWR.n4 VPWR.n3 5.012
R34 VPWR VPWR.n24 2.49
R35 VPWR.n23 VPWR.n22 0.231
R36 VPWR.n19 VPWR.n18 0.231
R37 VPWR.n16 VPWR.n15 0.231
R38 VPWR.n12 VPWR.n11 0.231
R39 VPWR.n9 VPWR.n8 0.231
R40 VPWR.n5 VPWR.n4 0.231
C0 VPWR a_230_351# 0.04fF
C1 B1 VPWR 0.03fF
C2 B1 a_230_351# 0.00fF
C3 A1 VPWR 0.09fF
C4 A1 a_230_351# 0.00fF
C5 B1 A1 0.04fF
C6 Y VPWR 0.16fF
C7 Y a_230_351# 0.08fF
C8 B1 Y 0.17fF
C9 Y A1 0.07fF
.ends

