magic
tech sky130A
magscale 1 2
timestamp 1678750074
<< nwell >>
rect -38 315 866 998
<< nmos >>
rect 195 47 225 223
rect 349 47 379 223
rect 503 47 533 223
rect 657 47 687 223
<< pmos >>
rect 195 351 225 913
rect 349 351 379 913
rect 503 351 533 913
rect 657 351 687 913
<< ndiff >>
rect 115 173 195 223
rect 115 139 138 173
rect 172 139 195 173
rect 115 105 195 139
rect 115 71 138 105
rect 172 71 195 105
rect 115 47 195 71
rect 225 105 349 223
rect 225 71 236 105
rect 270 71 304 105
rect 338 71 349 105
rect 225 47 349 71
rect 379 173 503 223
rect 379 139 424 173
rect 458 139 503 173
rect 379 105 503 139
rect 379 71 424 105
rect 458 71 503 105
rect 379 47 503 71
rect 533 215 657 223
rect 533 181 544 215
rect 578 181 612 215
rect 646 181 657 215
rect 533 47 657 181
rect 687 173 767 223
rect 687 139 710 173
rect 744 139 767 173
rect 687 105 767 139
rect 687 71 710 105
rect 744 71 767 105
rect 687 47 767 71
<< pdiff >>
rect 115 889 195 913
rect 115 855 138 889
rect 172 855 195 889
rect 115 821 195 855
rect 115 787 138 821
rect 172 787 195 821
rect 115 753 195 787
rect 115 719 138 753
rect 172 719 195 753
rect 115 685 195 719
rect 115 651 138 685
rect 172 651 195 685
rect 115 617 195 651
rect 115 583 138 617
rect 172 583 195 617
rect 115 549 195 583
rect 115 515 138 549
rect 172 515 195 549
rect 115 351 195 515
rect 225 351 349 913
rect 379 889 503 913
rect 379 855 425 889
rect 459 855 503 889
rect 379 821 503 855
rect 379 787 425 821
rect 459 787 503 821
rect 379 753 503 787
rect 379 719 425 753
rect 459 719 503 753
rect 379 685 503 719
rect 379 651 425 685
rect 459 651 503 685
rect 379 617 503 651
rect 379 583 425 617
rect 459 583 503 617
rect 379 549 503 583
rect 379 515 425 549
rect 459 515 503 549
rect 379 351 503 515
rect 533 351 657 913
rect 687 889 767 913
rect 687 855 710 889
rect 744 855 767 889
rect 687 821 767 855
rect 687 787 710 821
rect 744 787 767 821
rect 687 753 767 787
rect 687 719 710 753
rect 744 719 767 753
rect 687 685 767 719
rect 687 651 710 685
rect 744 651 767 685
rect 687 617 767 651
rect 687 583 710 617
rect 744 583 767 617
rect 687 549 767 583
rect 687 515 710 549
rect 744 515 767 549
rect 687 351 767 515
<< ndiffc >>
rect 138 139 172 173
rect 138 71 172 105
rect 236 71 270 105
rect 304 71 338 105
rect 424 139 458 173
rect 424 71 458 105
rect 544 181 578 215
rect 612 181 646 215
rect 710 139 744 173
rect 710 71 744 105
<< pdiffc >>
rect 138 855 172 889
rect 138 787 172 821
rect 138 719 172 753
rect 138 651 172 685
rect 138 583 172 617
rect 138 515 172 549
rect 425 855 459 889
rect 425 787 459 821
rect 425 719 459 753
rect 425 651 459 685
rect 425 583 459 617
rect 425 515 459 549
rect 710 855 744 889
rect 710 787 744 821
rect 710 719 744 753
rect 710 651 744 685
rect 710 583 744 617
rect 710 515 744 549
<< psubdiff >>
rect 36 173 115 223
rect 36 139 59 173
rect 93 139 115 173
rect 36 105 115 139
rect 36 71 59 105
rect 93 71 115 105
rect 36 47 115 71
<< nsubdiff >>
rect 36 889 115 913
rect 36 855 59 889
rect 93 855 115 889
rect 36 821 115 855
rect 36 787 59 821
rect 93 787 115 821
rect 36 753 115 787
rect 36 719 59 753
rect 93 719 115 753
rect 36 685 115 719
rect 36 651 59 685
rect 93 651 115 685
rect 36 617 115 651
rect 36 583 59 617
rect 93 583 115 617
rect 36 549 115 583
rect 36 515 59 549
rect 93 515 115 549
rect 36 351 115 515
<< psubdiffcont >>
rect 59 139 93 173
rect 59 71 93 105
<< nsubdiffcont >>
rect 59 855 93 889
rect 59 787 93 821
rect 59 719 93 753
rect 59 651 93 685
rect 59 583 93 617
rect 59 515 93 549
<< poly >>
rect 195 913 225 939
rect 349 913 379 939
rect 503 913 533 939
rect 657 913 687 939
rect 195 314 225 351
rect 349 314 379 351
rect 503 314 533 351
rect 657 314 687 351
rect 61 304 225 314
rect 61 270 77 304
rect 111 270 145 304
rect 179 270 225 304
rect 61 260 225 270
rect 267 304 401 314
rect 267 270 283 304
rect 317 270 351 304
rect 385 270 401 304
rect 267 260 401 270
rect 443 304 579 314
rect 443 270 459 304
rect 493 270 527 304
rect 561 270 579 304
rect 443 260 579 270
rect 657 304 797 314
rect 657 270 679 304
rect 713 270 747 304
rect 781 270 797 304
rect 657 260 797 270
rect 195 223 225 260
rect 349 223 379 260
rect 503 223 533 260
rect 657 223 687 260
rect 195 21 225 47
rect 349 21 379 47
rect 503 21 533 47
rect 657 21 687 47
<< polycont >>
rect 77 270 111 304
rect 145 270 179 304
rect 283 270 317 304
rect 351 270 385 304
rect 459 270 493 304
rect 527 270 561 304
rect 679 270 713 304
rect 747 270 781 304
<< locali >>
rect 0 943 29 977
rect 63 943 121 977
rect 155 943 213 977
rect 247 943 305 977
rect 339 943 397 977
rect 431 943 489 977
rect 523 943 581 977
rect 615 943 673 977
rect 707 943 765 977
rect 799 943 828 977
rect 59 889 172 943
rect 93 855 138 889
rect 59 821 172 855
rect 93 787 138 821
rect 59 753 172 787
rect 93 719 138 753
rect 59 685 172 719
rect 93 651 138 685
rect 59 617 172 651
rect 93 583 138 617
rect 59 549 172 583
rect 93 515 138 549
rect 59 499 172 515
rect 425 889 459 905
rect 425 821 459 855
rect 425 753 459 787
rect 425 685 459 719
rect 425 617 459 651
rect 425 549 459 583
rect 710 889 744 943
rect 710 821 744 855
rect 710 753 744 787
rect 710 685 744 719
rect 710 617 744 651
rect 710 549 744 583
rect 459 515 644 533
rect 425 499 644 515
rect 710 499 744 515
rect 77 304 179 406
rect 111 270 145 304
rect 77 254 179 270
rect 283 304 385 406
rect 317 270 351 304
rect 283 254 385 270
rect 459 304 561 406
rect 493 270 527 304
rect 459 254 561 270
rect 595 215 644 499
rect 679 304 781 406
rect 713 270 747 304
rect 679 254 781 270
rect 59 173 93 189
rect 59 105 93 139
rect 59 17 93 71
rect 138 173 459 189
rect 172 139 424 173
rect 458 139 459 173
rect 527 181 544 215
rect 578 181 612 215
rect 646 181 662 215
rect 527 147 662 181
rect 710 173 744 191
rect 138 105 172 139
rect 424 105 459 139
rect 138 51 172 71
rect 220 71 236 105
rect 270 71 304 105
rect 338 71 354 105
rect 220 17 354 71
rect 458 85 459 105
rect 710 105 744 139
rect 458 71 710 85
rect 424 51 744 71
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 943 63 977
rect 121 943 155 977
rect 213 943 247 977
rect 305 943 339 977
rect 397 943 431 977
rect 489 943 523 977
rect 581 943 615 977
rect 673 943 707 977
rect 765 943 799 977
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 977 828 1000
rect 0 943 29 977
rect 63 943 121 977
rect 155 943 213 977
rect 247 943 305 977
rect 339 943 397 977
rect 431 943 489 977
rect 523 943 581 977
rect 615 943 673 977
rect 707 943 765 977
rect 799 943 828 977
rect 0 920 828 943
rect 0 17 828 40
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -40 828 -17
<< labels >>
flabel locali s 121 343 155 377 0 FreeSans 240 0 0 0 A2
port 0 nsew signal input
flabel locali s 305 343 339 377 0 FreeSans 240 0 0 0 A1
port 1 nsew signal input
flabel locali s 489 343 523 377 0 FreeSans 240 0 0 0 B1
port 2 nsew signal input
flabel locali s 690 343 724 377 0 FreeSans 240 0 0 0 B2
port 3 nsew signal input
flabel metal1 s 397 943 431 977 0 FreeSans 240 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 397 -17 431 17 0 FreeSans 240 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 603 343 637 377 0 FreeSans 240 0 0 0 Y
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 960
string LEFclass CORE
string LEForigin 0 0
<< end >>
