* NGSPICE file created from thesis_oai22.ext - technology: sky130A

.subckt thesis_oai22 A2 A1 B1 B2 Y VPWR VGND
X0 Y.t0 A1.t0 a_225_351# VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.8711 pd=3.43 as=0.8711 ps=3.43 w=2.81 l=0.15
X1 a_115_47# A1.t1 VGND.t0 VGND sky130_fd_pr__nfet_01v8 ad=0.2728 pd=1.5 as=0.2728 ps=1.5 w=0.88 l=0.15
X2 Y.t1 B1.t0 a_115_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2728 pd=1.5 as=0.2728 ps=1.5 w=0.88 l=0.15
X3 a_533_351# B1.t1 Y.t2 VPWR.t1 sky130_fd_pr__pfet_01v8 ad=0.8711 pd=3.43 as=0.8711 ps=3.43 w=2.81 l=0.15
X4 VPWR.t3 B2.t0 a_533_351# VPWR.t2 sky130_fd_pr__pfet_01v8 ad=1.124 pd=6.42 as=0.8711 ps=3.43 w=2.81 l=0.15
X5 a_115_47# B2.t1 Y.t3 VGND sky130_fd_pr__nfet_01v8 ad=0.352 pd=2.56 as=0.2728 ps=1.5 w=0.88 l=0.15
X6 a_225_351# A2.t0 VPWR.t5 VPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.8711 pd=3.43 as=1.124 ps=6.42 w=2.81 l=0.15
X7 VGND.t1 A2.t1 a_115_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2728 pd=1.5 as=0.352 ps=2.56 w=0.88 l=0.15
R0 A1.n0 A1.t0 510.919
R1 A1.n0 A1.t1 200.832
R2 A1 A1.n0 51.894
R3 Y Y.n0 182.512
R4 Y Y.n1 73.413
R5 Y.n1 Y.t1 38.728
R6 Y.n1 Y.t3 37.012
R7 Y.n0 Y.t0 22.083
R8 Y.n0 Y.t2 21.382
R9 VPWR.t1 VPWR.t2 214.202
R10 VPWR.t0 VPWR.t1 214.202
R11 VPWR.t4 VPWR.t0 214.202
R12 VPWR.n14 VPWR.t4 186.383
R13 VPWR.n13 VPWR.n12 144.35
R14 VPWR.n17 VPWR.t3 131.688
R15 VPWR.n16 VPWR.n15 125.642
R16 VPWR.n6 VPWR.n5 92.5
R17 VPWR.n9 VPWR.n1 92.5
R18 VPWR.n7 VPWR.n2 92.5
R19 VPWR.n11 VPWR.n10 92.5
R20 VPWR.n1 VPWR.n0 33.142
R21 VPWR.n5 VPWR.n4 33.142
R22 VPWR.n15 VPWR.n14 29.68
R23 VPWR.n12 VPWR.t5 14.021
R24 VPWR.n17 VPWR.n16 13.143
R25 VPWR.n11 VPWR.n9 7.702
R26 VPWR.n7 VPWR.n6 7.702
R27 VPWR.n16 VPWR.n13 3.801
R28 VPWR.n8 VPWR.n7 3.801
R29 VPWR.n13 VPWR.n11 3.801
R30 VPWR.n9 VPWR.n8 3.801
R31 VPWR.n6 VPWR.n3 3.801
R32 VPWR.n17 VPWR 0.001
R33 VGND VGND.n0 39.652
R34 VGND.n0 VGND.t1 37.812
R35 VGND.n0 VGND.t0 37.611
R36 B1.n0 B1.t1 510.919
R37 B1.n0 B1.t0 200.832
R38 B1 B1.n0 54.473
R39 B2.n0 B2.t0 510.919
R40 B2.n0 B2.t1 200.832
R41 B2 B2.n0 71.483
R42 A2.n0 A2.t0 510.919
R43 A2.n0 A2.t1 200.832
R44 A2 A2.n0 93.395
C0 A1 B1 0.08fF
C1 A2 Y 0.00fF
C2 A2 a_225_351# 0.00fF
C3 A2 A1 0.07fF
C4 VPWR a_115_47# 0.04fF
C5 B2 a_533_351# 0.00fF
C6 Y B2 0.09fF
C7 B1 a_115_47# 0.04fF
C8 A2 a_115_47# 0.08fF
C9 VPWR B1 0.02fF
C10 a_115_47# B2 0.08fF
C11 Y a_533_351# 0.11fF
C12 A2 VPWR 0.09fF
C13 Y a_225_351# 0.02fF
C14 A1 Y 0.02fF
C15 A1 a_225_351# 0.04fF
C16 VPWR B2 0.13fF
C17 B1 B2 0.03fF
C18 a_115_47# Y 0.13fF
C19 a_115_47# a_225_351# 0.02fF
C20 A1 a_115_47# 0.08fF
C21 VPWR a_533_351# 0.05fF
C22 VPWR Y 0.19fF
C23 VPWR a_225_351# 0.05fF
C24 VPWR A1 0.03fF
C25 B1 a_533_351# 0.01fF
C26 B1 Y 0.16fF
.ends

