* NGSPICE file created from thesis_aoi211.ext - technology: sky130A

.subckt thesis_aoi211 A2 A1 B1 C1 Y VPWR VGND
X0 a_115_351# A1.t0 VPWR.t1 VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.8711 pd=3.43 as=0.8711 ps=3.43 w=2.81 l=0.15
X1 Y.t0 A1.t1 a_225_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2728 pd=1.5 as=0.2728 ps=1.5 w=0.88 l=0.15
X2 VGND.t0 B1.t0 Y.t1 VGND sky130_fd_pr__nfet_01v8 ad=0.2728 pd=1.5 as=0.2728 ps=1.5 w=0.88 l=0.15
X3 a_533_351# B1.t1 a_115_351# VPWR.t2 sky130_fd_pr__pfet_01v8 ad=0.8711 pd=3.43 as=0.8711 ps=3.43 w=2.81 l=0.15
X4 Y.t2 C1.t0 a_533_351# VPWR.t3 sky130_fd_pr__pfet_01v8 ad=1.124 pd=6.42 as=0.8711 ps=3.43 w=2.81 l=0.15
X5 Y.t3 C1.t1 VGND.t2 VGND sky130_fd_pr__nfet_01v8 ad=0.352 pd=2.56 as=0.2728 ps=1.5 w=0.88 l=0.15
X6 VPWR.t5 A2.t0 a_115_351# VPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.8711 pd=3.43 as=1.124 ps=6.42 w=2.81 l=0.15
X7 a_225_47# A2.t1 VGND.t1 VGND sky130_fd_pr__nfet_01v8 ad=0.2728 pd=1.5 as=0.352 ps=2.56 w=0.88 l=0.15
R0 A1.n0 A1.t0 510.919
R1 A1.n0 A1.t1 200.832
R2 A1 A1.n0 52.258
R3 VPWR.n1 VPWR.t4 280.503
R4 VPWR.t2 VPWR.t3 214.202
R5 VPWR.t0 VPWR.t2 214.202
R6 VPWR.t4 VPWR.t0 214.202
R7 VPWR.n1 VPWR.n0 43.925
R8 VPWR.n0 VPWR.t1 19.394
R9 VPWR.n0 VPWR.t5 19.394
R10 VPWR VPWR.n1 0.239
R11 Y.n2 Y.n1 158.062
R12 Y.n1 Y.t3 124.966
R13 Y.n1 Y.n0 118.174
R14 Y.n2 Y.t2 62.833
R15 Y.n0 Y.t1 42.272
R16 Y.n0 Y.t0 42.272
R17 Y Y.n2 10.386
R18 VGND.n3 VGND.n2 94.773
R19 VGND.n1 VGND.n0 92.5
R20 VGND.n8 VGND.t1 86.992
R21 VGND.n2 VGND.t2 19.09
R22 VGND.n0 VGND.t0 19.09
R23 VGND.n5 VGND.n4 4.65
R24 VGND.n7 VGND.n6 4.65
R25 VGND.n3 VGND.n1 4.459
R26 VGND.n5 VGND.n3 3.392
R27 VGND VGND.n8 0.197
R28 VGND.n7 VGND.n5 0.143
R29 VGND VGND.n7 0.026
R30 B1.n0 B1.t1 510.919
R31 B1.n0 B1.t0 200.832
R32 B1 B1.n0 54.744
R33 C1.n0 C1.t0 510.919
R34 C1.n0 C1.t1 200.832
R35 C1 C1.n0 71.721
R36 A2.n0 A2.t0 510.919
R37 A2.n0 A2.t1 200.832
R38 A2 A2.n0 93.698
C0 B1 a_533_351# 0.01fF
C1 C1 a_533_351# 0.00fF
C2 a_115_351# a_533_351# 0.03fF
C3 a_225_47# a_115_351# 0.02fF
C4 a_225_47# A1 0.02fF
C5 Y a_533_351# 0.10fF
C6 a_225_47# Y 0.01fF
C7 VPWR a_533_351# 0.04fF
C8 B1 C1 0.03fF
C9 a_115_351# B1 0.04fF
C10 a_115_351# C1 0.00fF
C11 A2 a_115_351# 0.09fF
C12 a_225_47# VPWR 0.00fF
C13 B1 A1 0.07fF
C14 a_115_351# A1 0.10fF
C15 A2 A1 0.07fF
C16 B1 Y 0.14fF
C17 Y C1 0.23fF
C18 a_115_351# Y 0.07fF
C19 A2 Y 0.00fF
C20 Y A1 0.01fF
C21 B1 VPWR 0.02fF
C22 VPWR C1 0.03fF
C23 a_115_351# VPWR 0.70fF
C24 A2 VPWR 0.06fF
C25 VPWR A1 0.05fF
C26 VPWR Y 0.11fF
.ends

