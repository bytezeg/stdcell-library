VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO thesis_aoi211
  CLASS CORE ;
  FOREIGN thesis_aoi211 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 4.800 ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.553500 ;
    PORT
      LAYER li1 ;
        RECT 0.385 1.270 0.895 1.915 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.553500 ;
    PORT
      LAYER li1 ;
        RECT 1.415 1.270 1.925 1.915 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.553500 ;
    PORT
      LAYER li1 ;
        RECT 2.295 1.270 2.805 1.915 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.553500 ;
    PORT
      LAYER li1 ;
        RECT 3.390 1.270 3.905 1.915 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.021600 ;
    PORT
      LAYER li1 ;
        RECT 3.550 3.650 3.720 4.535 ;
        RECT 3.550 2.335 3.725 3.650 ;
        RECT 2.975 2.165 3.725 2.335 ;
        RECT 2.975 1.005 3.145 2.165 ;
        RECT 2.120 0.830 3.720 1.005 ;
        RECT 2.120 0.255 2.290 0.830 ;
        RECT 3.550 0.255 3.720 0.830 ;
    END
  END Y
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.575 4.330 4.990 ;
      LAYER li1 ;
        RECT 0.000 4.715 4.140 4.885 ;
        RECT 0.295 2.155 0.465 4.715 ;
        RECT 1.180 2.495 1.695 4.715 ;
      LAYER mcon ;
        RECT 0.140 4.715 0.310 4.885 ;
        RECT 0.605 4.715 0.775 4.885 ;
        RECT 1.065 4.715 1.235 4.885 ;
        RECT 1.525 4.715 1.695 4.885 ;
        RECT 1.985 4.715 2.155 4.885 ;
        RECT 2.445 4.715 2.615 4.885 ;
        RECT 2.905 4.715 3.075 4.885 ;
        RECT 3.365 4.715 3.535 4.885 ;
        RECT 3.825 4.715 3.995 4.885 ;
      LAYER met1 ;
        RECT 0.000 4.600 4.140 5.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.290 0.085 0.920 0.950 ;
        RECT 2.635 0.085 3.310 0.525 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.200 4.140 0.200 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.690 2.325 0.860 4.545 ;
        RECT 2.120 2.325 2.290 4.545 ;
        RECT 0.690 2.155 2.290 2.325 ;
  END
END thesis_aoi211
END LIBRARY

