* NGSPICE file created from thesis_inv.ext - technology: sky130A

.subckt inverter VPWR Y A VGND
X0 Y.t1 A.t0 VPWR.t1 VPWR.t0 sky130_fd_pr__pfet_01v8 ad=1.25045 pd=6.51 as=1.2364 ps=6.5 w=2.81 l=0.15
X1 Y.t0 A.t1 VGND.t0 VGND sky130_fd_pr__nfet_01v8 ad=0.3916 pd=2.65 as=0.3872 ps=2.64 w=0.88 l=0.15
R0 A.n0 A.t0 510.919
R1 A.n0 A.t1 200.832
R2 A A.n0 93.033
R3 VPWR.n14 VPWR.t0 205.555
R4 VPWR.n13 VPWR.n12 144.503
R5 VPWR.n16 VPWR.n15 123.152
R6 VPWR.n6 VPWR.n5 92.5
R7 VPWR.n9 VPWR.n1 92.5
R8 VPWR.n7 VPWR.n2 92.5
R9 VPWR.n11 VPWR.n10 92.5
R10 VPWR.n15 VPWR.n14 30.925
R11 VPWR.n1 VPWR.n0 30.652
R12 VPWR.n5 VPWR.n4 30.652
R13 VPWR.n12 VPWR.t1 15.423
R14 VPWR VPWR.n16 10.137
R15 VPWR.n11 VPWR.n9 7.076
R16 VPWR.n7 VPWR.n6 7.076
R17 VPWR.n16 VPWR.n13 3.496
R18 VPWR.n8 VPWR.n7 3.496
R19 VPWR.n13 VPWR.n11 3.496
R20 VPWR.n9 VPWR.n8 3.496
R21 VPWR.n6 VPWR.n3 3.496
R22 Y Y.t0 116.091
R23 Y Y.t1 58.49
R24 VGND VGND.t0 87.219
C0 VPWR A 0.13fF
C1 Y A 0.11fF
C2 Y VPWR 0.22fF
.ends

