* NGSPICE file created from thesis_oai211.ext - technology: sky130A

.subckt thesis_oai211 A2 A1 B1 C1 Y VPWR VGND
X0 Y.t0 A1.t0 a_225_351# VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.8711 pd=3.43 as=0.8711 ps=3.43 w=2.81 l=0.15
X1 a_115_47# A1.t1 VGND.t0 VGND sky130_fd_pr__nfet_01v8 ad=0.2728 pd=1.5 as=0.2728 ps=1.5 w=0.88 l=0.15
X2 a_533_47# B1.t0 a_115_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2728 pd=1.5 as=0.2728 ps=1.5 w=0.88 l=0.15
X3 VPWR.t2 B1.t1 Y.t1 VPWR.t1 sky130_fd_pr__pfet_01v8 ad=0.8711 pd=3.43 as=0.8711 ps=3.43 w=2.81 l=0.15
X4 Y.t2 C1.t0 VPWR.t4 VPWR.t3 sky130_fd_pr__pfet_01v8 ad=1.124 pd=6.42 as=0.8711 ps=3.43 w=2.81 l=0.15
X5 Y.t3 C1.t1 a_533_47# VGND sky130_fd_pr__nfet_01v8 ad=0.352 pd=2.56 as=0.2728 ps=1.5 w=0.88 l=0.15
X6 a_225_351# A2.t0 VPWR.t6 VPWR.t5 sky130_fd_pr__pfet_01v8 ad=0.8711 pd=3.43 as=1.124 ps=6.42 w=2.81 l=0.15
X7 VGND.t1 A2.t1 a_115_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2728 pd=1.5 as=0.352 ps=2.56 w=0.88 l=0.15
R0 A1.n0 A1.t0 510.919
R1 A1.n0 A1.t1 200.832
R2 A1 A1.n0 52.203
R3 Y Y.t3 149.921
R4 Y.n1 Y.n0 118.066
R5 Y.n1 Y.t2 117.495
R6 Y Y.n1 63.247
R7 Y.n0 Y.t1 22.083
R8 Y.n0 Y.t0 21.382
R9 VPWR.t1 VPWR.t3 214.202
R10 VPWR.t0 VPWR.t1 214.202
R11 VPWR.t5 VPWR.t0 214.202
R12 VPWR.n17 VPWR.t5 186.383
R13 VPWR.n16 VPWR.n15 144.35
R14 VPWR.n19 VPWR.n18 125.642
R15 VPWR.n6 VPWR.n5 96.302
R16 VPWR.n8 VPWR.n7 92.5
R17 VPWR.n12 VPWR.n1 92.5
R18 VPWR.n11 VPWR.n2 92.5
R19 VPWR.n9 VPWR.n4 92.5
R20 VPWR.n14 VPWR.n13 92.5
R21 VPWR.n21 VPWR.n20 47.854
R22 VPWR.n1 VPWR.n0 33.142
R23 VPWR.n4 VPWR.n3 33.142
R24 VPWR.n18 VPWR.n17 29.68
R25 VPWR.n20 VPWR.t2 19.718
R26 VPWR.n20 VPWR.t4 19.718
R27 VPWR.n15 VPWR.t6 14.021
R28 VPWR.n21 VPWR.n19 13.142
R29 VPWR.n14 VPWR.n12 7.702
R30 VPWR.n12 VPWR.n11 7.702
R31 VPWR.n9 VPWR.n8 7.702
R32 VPWR.n19 VPWR.n16 3.801
R33 VPWR.n10 VPWR.n9 3.801
R34 VPWR.n16 VPWR.n14 3.801
R35 VPWR.n11 VPWR.n10 3.801
R36 VPWR.n8 VPWR.n6 3.801
R37 VPWR VPWR.n21 0.001
R38 VGND VGND.n0 39.652
R39 VGND.n0 VGND.t1 37.812
R40 VGND.n0 VGND.t0 37.611
R41 B1.n0 B1.t1 510.919
R42 B1.n0 B1.t0 200.832
R43 B1 B1.n0 54.703
R44 C1.n0 C1.t0 510.919
R45 C1.n0 C1.t1 200.832
R46 C1 C1.n0 66.471
R47 A2.n0 A2.t0 510.919
R48 A2.n0 A2.t1 200.832
R49 A2 A2.n0 93.652
C0 A1 A2 0.07fF
C1 a_533_47# B1 0.01fF
C2 VPWR A2 0.10fF
C3 C1 Y 0.22fF
C4 a_115_47# C1 0.00fF
C5 a_115_47# Y 0.04fF
C6 A1 B1 0.07fF
C7 a_225_351# Y 0.02fF
C8 VPWR B1 0.03fF
C9 a_115_47# a_225_351# 0.02fF
C10 a_533_47# Y 0.03fF
C11 a_533_47# a_115_47# 0.00fF
C12 A1 Y 0.01fF
C13 C1 VPWR 0.04fF
C14 VPWR Y 0.53fF
C15 A1 a_115_47# 0.08fF
C16 a_115_47# VPWR 0.04fF
C17 A1 a_225_351# 0.04fF
C18 a_225_351# VPWR 0.05fF
C19 A2 Y 0.00fF
C20 a_533_47# VPWR 0.00fF
C21 a_115_47# A2 0.08fF
C22 a_225_351# A2 0.00fF
C23 C1 B1 0.03fF
C24 Y B1 0.15fF
C25 A1 VPWR 0.03fF
C26 a_115_47# B1 0.01fF
.ends

