magic
tech sky130A
magscale 1 2
timestamp 1678764467
<< nwell >>
rect -38 315 682 998
<< nmos >>
rect 186 47 216 223
rect 325 47 355 223
rect 464 47 494 223
<< pmos >>
rect 186 351 216 913
rect 325 351 355 913
rect 464 351 494 913
<< ndiff >>
rect 111 173 186 223
rect 111 139 132 173
rect 166 139 186 173
rect 111 105 186 139
rect 111 71 132 105
rect 166 71 186 105
rect 111 47 186 71
rect 216 157 325 223
rect 216 123 253 157
rect 287 123 325 157
rect 216 89 325 123
rect 216 55 253 89
rect 287 55 325 89
rect 216 47 325 55
rect 355 169 464 223
rect 355 135 393 169
rect 427 135 464 169
rect 355 101 464 135
rect 355 67 393 101
rect 427 67 464 101
rect 355 47 464 67
rect 494 169 569 223
rect 494 135 514 169
rect 548 135 569 169
rect 494 101 569 135
rect 494 67 514 101
rect 548 67 569 101
rect 494 47 569 67
<< pdiff >>
rect 111 889 186 913
rect 111 855 141 889
rect 175 855 186 889
rect 111 821 186 855
rect 111 787 141 821
rect 175 787 186 821
rect 111 753 186 787
rect 111 719 141 753
rect 175 719 186 753
rect 111 685 186 719
rect 111 651 141 685
rect 175 651 186 685
rect 111 617 186 651
rect 111 583 141 617
rect 175 583 186 617
rect 111 351 186 583
rect 216 351 325 913
rect 355 889 464 913
rect 355 855 392 889
rect 426 855 464 889
rect 355 821 464 855
rect 355 787 392 821
rect 426 787 464 821
rect 355 753 464 787
rect 355 719 392 753
rect 426 719 464 753
rect 355 685 464 719
rect 355 651 392 685
rect 426 651 464 685
rect 355 617 464 651
rect 355 583 392 617
rect 426 583 464 617
rect 355 351 464 583
rect 494 889 569 913
rect 494 855 515 889
rect 549 855 569 889
rect 494 821 569 855
rect 494 787 515 821
rect 549 787 569 821
rect 494 753 569 787
rect 494 719 515 753
rect 549 719 569 753
rect 494 685 569 719
rect 494 651 515 685
rect 549 651 569 685
rect 494 617 569 651
rect 494 583 515 617
rect 549 583 569 617
rect 494 351 569 583
<< ndiffc >>
rect 132 139 166 173
rect 132 71 166 105
rect 253 123 287 157
rect 253 55 287 89
rect 393 135 427 169
rect 393 67 427 101
rect 514 135 548 169
rect 514 67 548 101
<< pdiffc >>
rect 141 855 175 889
rect 141 787 175 821
rect 141 719 175 753
rect 141 651 175 685
rect 141 583 175 617
rect 392 855 426 889
rect 392 787 426 821
rect 392 719 426 753
rect 392 651 426 685
rect 392 583 426 617
rect 515 855 549 889
rect 515 787 549 821
rect 515 719 549 753
rect 515 651 549 685
rect 515 583 549 617
<< psubdiff >>
rect 36 173 111 223
rect 36 139 56 173
rect 90 139 111 173
rect 36 105 111 139
rect 36 71 56 105
rect 90 71 111 105
rect 36 47 111 71
<< nsubdiff >>
rect 36 889 111 913
rect 36 855 53 889
rect 87 855 111 889
rect 36 821 111 855
rect 36 787 53 821
rect 87 787 111 821
rect 36 753 111 787
rect 36 719 53 753
rect 87 719 111 753
rect 36 685 111 719
rect 36 651 53 685
rect 87 651 111 685
rect 36 617 111 651
rect 36 583 53 617
rect 87 583 111 617
rect 36 351 111 583
<< psubdiffcont >>
rect 56 139 90 173
rect 56 71 90 105
<< nsubdiffcont >>
rect 53 855 87 889
rect 53 787 87 821
rect 53 719 87 753
rect 53 651 87 685
rect 53 583 87 617
<< poly >>
rect 186 913 216 939
rect 325 913 355 939
rect 464 913 494 939
rect 186 314 216 351
rect 325 314 355 351
rect 464 314 494 351
rect 52 304 216 314
rect 52 270 68 304
rect 102 270 136 304
rect 170 270 216 304
rect 52 260 216 270
rect 258 304 394 314
rect 258 270 276 304
rect 310 270 344 304
rect 378 270 394 304
rect 258 260 394 270
rect 436 304 572 314
rect 436 270 452 304
rect 486 270 520 304
rect 554 270 572 304
rect 186 223 216 260
rect 325 223 355 260
rect 436 259 572 270
rect 464 223 494 259
rect 186 21 216 47
rect 325 21 355 47
rect 464 21 494 47
<< polycont >>
rect 68 270 102 304
rect 136 270 170 304
rect 276 270 310 304
rect 344 270 378 304
rect 452 270 486 304
rect 520 270 554 304
<< locali >>
rect 0 943 29 977
rect 63 943 121 977
rect 155 943 213 977
rect 247 943 305 977
rect 339 943 397 977
rect 431 943 489 977
rect 523 943 581 977
rect 615 943 644 977
rect 53 889 175 943
rect 87 855 141 889
rect 53 821 175 855
rect 87 787 141 821
rect 53 753 175 787
rect 87 719 141 753
rect 53 685 175 719
rect 87 651 141 685
rect 53 617 175 651
rect 87 583 141 617
rect 53 565 175 583
rect 392 889 426 909
rect 392 821 426 855
rect 392 753 426 787
rect 392 685 426 719
rect 392 617 426 651
rect 392 473 426 583
rect 515 889 549 943
rect 515 821 549 855
rect 515 753 549 787
rect 515 685 549 719
rect 515 617 549 651
rect 515 565 549 583
rect 392 437 640 473
rect 52 304 186 403
rect 52 270 68 304
rect 102 270 136 304
rect 170 270 186 304
rect 260 304 394 403
rect 260 270 276 304
rect 310 270 344 304
rect 378 270 394 304
rect 436 304 572 403
rect 436 270 452 304
rect 486 270 520 304
rect 554 270 572 304
rect 606 236 640 437
rect 132 191 427 225
rect 56 173 90 189
rect 56 105 90 139
rect 56 17 90 71
rect 132 173 166 191
rect 393 169 427 191
rect 132 105 166 139
rect 132 51 166 71
rect 237 123 253 157
rect 287 123 303 157
rect 237 89 303 123
rect 237 55 253 89
rect 287 55 303 89
rect 237 17 303 55
rect 393 101 427 135
rect 393 51 427 67
rect 514 202 640 236
rect 514 169 548 202
rect 514 101 548 135
rect 514 51 548 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 943 63 977
rect 121 943 155 977
rect 213 943 247 977
rect 305 943 339 977
rect 397 943 431 977
rect 489 943 523 977
rect 581 943 615 977
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 977 644 1000
rect 0 943 29 977
rect 63 943 121 977
rect 155 943 213 977
rect 247 943 305 977
rect 339 943 397 977
rect 431 943 489 977
rect 523 943 581 977
rect 615 943 644 977
rect 0 920 644 943
rect 0 17 644 40
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -40 644 -17
<< labels >>
flabel metal1 s 305 -17 339 17 0 FreeSans 240 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 110 343 144 377 0 FreeSans 240 0 0 0 A1
port 0 nsew signal input
flabel locali s 294 343 328 377 0 FreeSans 240 0 0 0 A2
port 1 nsew signal input
flabel locali s 476 343 510 377 0 FreeSans 240 0 0 0 B1
port 2 nsew signal input
flabel locali s 606 343 640 377 0 FreeSans 240 0 0 0 Y
port 3 nsew signal output
flabel metal1 s 305 943 339 977 0 FreeSans 240 0 0 0 VPWR
port 4 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 644 960
string LEFclass CORE
string LEForigin 0 0
<< end >>
