* NGSPICE file created from thesis_nand2.ext - technology: sky130A

.subckt thesis_nand2 A1 B1 Y VPWR VGND
X0 Y.t2 B1.t0 a_230_47# VGND sky130_fd_pr__nfet_01v8 ad=0.3608 pd=2.58 as=0.1804 ps=1.29 w=0.88 l=0.15
X1 a_230_47# A1.t0 VGND.t0 VGND sky130_fd_pr__nfet_01v8 ad=0.1804 pd=1.29 as=0.3608 ps=2.58 w=0.88 l=0.15
X2 VPWR.t3 B1.t1 Y.t1 VPWR.t2 sky130_fd_pr__pfet_01v8 ad=1.1521 pd=6.44 as=0.57605 ps=3.22 w=2.81 l=0.15
X3 Y.t0 A1.t1 VPWR.t1 VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.57605 pd=3.22 as=1.2645 ps=6.52 w=2.81 l=0.15
R0 B1.n0 B1.t1 510.919
R1 B1.n0 B1.t0 200.832
R2 B1 B1.n0 52.922
R3 Y Y.t2 178.957
R4 Y Y.n0 111.431
R5 Y.n0 Y.t0 14.722
R6 Y.n0 Y.t1 14.021
R7 VGND VGND.t0 88.74
R8 A1.n0 A1.t1 510.919
R9 A1.n0 A1.t0 200.832
R10 A1 A1.n0 70.693
R11 VPWR.n24 VPWR.n1 292.5
R12 VPWR.n21 VPWR.t0 203.074
R13 VPWR.t0 VPWR.t2 155.783
R14 VPWR.n0 VPWR.t3 127.696
R15 VPWR.n23 VPWR.n22 127.045
R16 VPWR.n4 VPWR.n3 92.731
R17 VPWR.n5 VPWR.n2 92.5
R18 VPWR.n16 VPWR.n15 92.5
R19 VPWR.n12 VPWR.n11 92.5
R20 VPWR.n9 VPWR.n8 92.5
R21 VPWR.n19 VPWR.n18 92.5
R22 VPWR.n15 VPWR.n14 34.545
R23 VPWR.n8 VPWR.n7 34.545
R24 VPWR.n22 VPWR.n21 28.978
R25 VPWR.n1 VPWR.t1 12.619
R26 VPWR.n25 VPWR.n24 6.554
R27 VPWR.n23 VPWR.n20 5.012
R28 VPWR.n19 VPWR.n17 5.012
R29 VPWR.n16 VPWR.n13 5.012
R30 VPWR.n12 VPWR.n10 5.012
R31 VPWR.n9 VPWR.n6 5.012
R32 VPWR.n5 VPWR.n4 5.012
R33 VPWR VPWR.n25 2.49
R34 VPWR.n24 VPWR.n23 0.231
R35 VPWR.n20 VPWR.n19 0.231
R36 VPWR.n17 VPWR.n16 0.231
R37 VPWR.n13 VPWR.n12 0.231
R38 VPWR.n10 VPWR.n9 0.231
R39 VPWR.n6 VPWR.n5 0.231
R40 VPWR VPWR.n0 0.215
C0 Y VPWR 0.39fF
C1 Y a_230_47# 0.03fF
C2 B1 Y 0.16fF
C3 Y A1 0.08fF
C4 VPWR a_230_47# 0.00fF
C5 B1 VPWR 0.08fF
C6 A1 VPWR 0.09fF
C7 B1 A1 0.04fF
.ends

