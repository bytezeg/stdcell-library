magic
tech sky130A
magscale 1 2
timestamp 1682107102
<< nwell >>
rect -38 315 498 998
<< nmos >>
rect 200 47 230 223
rect 312 47 342 223
<< pmos >>
rect 200 351 230 913
rect 312 351 342 913
<< ndiff >>
rect 118 170 200 223
rect 118 136 138 170
rect 172 136 200 170
rect 118 102 200 136
rect 118 68 138 102
rect 172 68 200 102
rect 118 47 200 68
rect 230 157 312 223
rect 230 123 254 157
rect 288 123 312 157
rect 230 89 312 123
rect 230 55 254 89
rect 288 55 312 89
rect 230 47 312 55
rect 342 170 424 223
rect 342 136 366 170
rect 400 136 424 170
rect 342 102 424 136
rect 342 68 366 102
rect 400 68 424 102
rect 342 47 424 68
<< pdiff >>
rect 110 892 200 913
rect 110 858 147 892
rect 181 858 200 892
rect 110 824 200 858
rect 110 790 147 824
rect 181 790 200 824
rect 110 756 200 790
rect 110 722 147 756
rect 181 722 200 756
rect 110 688 200 722
rect 110 654 147 688
rect 181 654 200 688
rect 110 620 200 654
rect 110 586 147 620
rect 181 586 200 620
rect 110 351 200 586
rect 230 892 312 913
rect 230 858 255 892
rect 289 858 312 892
rect 230 824 312 858
rect 230 790 255 824
rect 289 790 312 824
rect 230 756 312 790
rect 230 722 255 756
rect 289 722 312 756
rect 230 688 312 722
rect 230 654 255 688
rect 289 654 312 688
rect 230 620 312 654
rect 230 586 255 620
rect 289 586 312 620
rect 230 351 312 586
rect 342 892 424 913
rect 342 858 366 892
rect 400 858 424 892
rect 342 824 424 858
rect 342 790 366 824
rect 400 790 424 824
rect 342 756 424 790
rect 342 722 366 756
rect 400 722 424 756
rect 342 688 424 722
rect 342 654 366 688
rect 400 654 424 688
rect 342 620 424 654
rect 342 586 366 620
rect 400 586 424 620
rect 342 552 424 586
rect 342 518 366 552
rect 400 518 424 552
rect 342 484 424 518
rect 342 450 366 484
rect 400 450 424 484
rect 342 351 424 450
<< ndiffc >>
rect 138 136 172 170
rect 138 68 172 102
rect 254 123 288 157
rect 254 55 288 89
rect 366 136 400 170
rect 366 68 400 102
<< pdiffc >>
rect 147 858 181 892
rect 147 790 181 824
rect 147 722 181 756
rect 147 654 181 688
rect 147 586 181 620
rect 255 858 289 892
rect 255 790 289 824
rect 255 722 289 756
rect 255 654 289 688
rect 255 586 289 620
rect 366 858 400 892
rect 366 790 400 824
rect 366 722 400 756
rect 366 654 400 688
rect 366 586 400 620
rect 366 518 400 552
rect 366 450 400 484
<< psubdiff >>
rect 36 173 118 223
rect 36 139 56 173
rect 90 139 118 173
rect 36 105 118 139
rect 36 71 56 105
rect 90 71 118 105
rect 36 47 118 71
<< nsubdiff >>
rect 36 889 110 913
rect 36 855 52 889
rect 86 855 110 889
rect 36 821 110 855
rect 36 787 52 821
rect 86 787 110 821
rect 36 753 110 787
rect 36 719 52 753
rect 86 719 110 753
rect 36 685 110 719
rect 36 651 52 685
rect 86 651 110 685
rect 36 617 110 651
rect 36 583 52 617
rect 86 583 110 617
rect 36 351 110 583
<< psubdiffcont >>
rect 56 139 90 173
rect 56 71 90 105
<< nsubdiffcont >>
rect 52 855 86 889
rect 52 787 86 821
rect 52 719 86 753
rect 52 651 86 685
rect 52 583 86 617
<< poly >>
rect 200 913 230 939
rect 312 913 342 939
rect 200 314 230 351
rect 312 314 342 351
rect 80 304 230 314
rect 80 270 109 304
rect 143 270 177 304
rect 211 270 230 304
rect 80 260 230 270
rect 272 304 407 314
rect 272 270 288 304
rect 322 270 356 304
rect 390 270 407 304
rect 272 260 407 270
rect 200 223 230 260
rect 312 223 342 260
rect 200 21 230 47
rect 312 21 342 47
<< polycont >>
rect 109 270 143 304
rect 177 270 211 304
rect 288 270 322 304
rect 356 270 390 304
<< locali >>
rect 0 943 29 977
rect 63 943 121 977
rect 155 943 213 977
rect 247 943 305 977
rect 339 943 397 977
rect 431 943 460 977
rect 36 889 100 943
rect 36 855 52 889
rect 86 855 100 889
rect 36 821 100 855
rect 36 787 52 821
rect 86 787 100 821
rect 36 753 100 787
rect 36 719 52 753
rect 86 719 100 753
rect 36 685 100 719
rect 36 651 52 685
rect 86 651 100 685
rect 36 617 100 651
rect 36 583 52 617
rect 86 583 100 617
rect 36 567 100 583
rect 135 892 202 908
rect 135 858 147 892
rect 181 858 202 892
rect 135 824 202 858
rect 135 790 147 824
rect 181 790 202 824
rect 135 756 202 790
rect 135 722 147 756
rect 181 722 202 756
rect 135 688 202 722
rect 135 654 147 688
rect 181 654 202 688
rect 135 620 202 654
rect 135 586 147 620
rect 181 586 202 620
rect 239 892 305 943
rect 239 858 255 892
rect 289 858 305 892
rect 239 824 305 858
rect 239 790 255 824
rect 289 790 305 824
rect 239 756 305 790
rect 239 722 255 756
rect 289 722 305 756
rect 239 688 305 722
rect 239 654 255 688
rect 289 654 305 688
rect 239 620 305 654
rect 239 586 255 620
rect 289 586 305 620
rect 366 892 400 908
rect 366 824 400 858
rect 366 756 400 790
rect 366 688 400 722
rect 366 620 400 654
rect 135 535 202 586
rect 366 552 400 586
rect 135 495 295 535
rect 93 304 227 432
rect 93 270 109 304
rect 143 270 177 304
rect 211 270 227 304
rect 261 320 295 495
rect 366 493 400 518
rect 366 484 459 493
rect 400 450 459 484
rect 366 433 459 450
rect 261 304 390 320
rect 261 270 288 304
rect 322 270 356 304
rect 261 254 390 270
rect 261 225 295 254
rect 134 191 295 225
rect 424 192 459 433
rect 36 173 100 189
rect 36 139 56 173
rect 90 139 100 173
rect 36 105 100 139
rect 36 71 56 105
rect 90 71 100 105
rect 36 17 100 71
rect 134 170 172 191
rect 134 136 138 170
rect 365 170 459 192
rect 134 102 172 136
rect 134 68 138 102
rect 134 52 172 68
rect 235 123 254 157
rect 288 123 309 157
rect 235 89 309 123
rect 235 55 254 89
rect 288 55 309 89
rect 235 17 309 55
rect 365 136 366 170
rect 400 158 459 170
rect 365 102 400 136
rect 365 68 366 102
rect 365 51 400 68
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 943 63 977
rect 121 943 155 977
rect 213 943 247 977
rect 305 943 339 977
rect 397 943 431 977
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 977 460 1000
rect 0 943 29 977
rect 63 943 121 977
rect 155 943 213 977
rect 247 943 305 977
rect 339 943 397 977
rect 431 943 460 977
rect 0 920 460 943
rect 0 17 460 40
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -40 460 -17
<< comment >>
rect 227 270 261 304
rect 160 220 194 254
rect 254 157 288 191
<< labels >>
flabel locali s 121 343 155 377 0 FreeSans 240 0 0 0 A1
port 0 nsew signal input
flabel metal1 s 121 943 155 977 0 FreeSans 240 0 0 0 VPWR
port 2 nsew
flabel metal1 s 213 -17 247 17 0 FreeSans 240 0 0 0 VGND
port 3 nsew
flabel locali s 425 274 459 308 0 FreeSans 240 0 0 0 Y
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 460 960
string LEFclass CORE
string LEForigin 0 0
<< end >>
