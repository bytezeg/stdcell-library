* NGSPICE file created from thesis_aoi21.ext - technology: sky130A

.subckt thesis_aoi21 A1 A2 B1 Y VPWR VGND
X0 VPWR.t4 A1.t0 a_116_351# VPWR.t3 sky130_fd_pr__pfet_01v8 ad=0.765725 pd=3.355 as=1.13805 ps=6.43 w=2.81 l=0.15
X1 Y.t0 A2.t0 a_227_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2398 pd=1.425 as=0.2398 ps=1.425 w=0.88 l=0.15
X2 Y.t1 B1.t0 a_116_351# VPWR.t2 sky130_fd_pr__pfet_01v8 ad=1.13805 pd=6.43 as=0.765725 ps=3.355 w=2.81 l=0.15
X3 VGND.t0 B1.t1 Y.t2 VGND sky130_fd_pr__nfet_01v8 ad=0.355875 pd=2.57 as=0.2398 ps=1.425 w=0.88 l=0.15
X4 a_227_47# A1.t1 VGND.t1 VGND sky130_fd_pr__nfet_01v8 ad=0.2398 pd=1.425 as=0.3564 ps=2.57 w=0.88 l=0.15
X5 a_116_351# A2.t1 VPWR.t1 VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.765725 pd=3.355 as=0.765725 ps=3.355 w=2.81 l=0.15
R0 A1.n0 A1.t0 510.919
R1 A1.n0 A1.t1 200.832
R2 A1 A1.n0 93.476
R3 VPWR.n1 VPWR.t3 287.357
R4 VPWR.t0 VPWR.t2 193.338
R5 VPWR.t3 VPWR.t0 193.338
R6 VPWR.n1 VPWR.n0 94.135
R7 VPWR.n0 VPWR.t4 19.279
R8 VPWR.n0 VPWR.t1 18.928
R9 VPWR VPWR.n1 0.116
R10 A2.n0 A2.t1 510.919
R11 A2.n0 A2.t0 200.832
R12 A2 A2.n0 54.282
R13 Y.n2 Y.n1 265.458
R14 Y.n2 Y.n0 87.113
R15 Y.n1 Y.t0 37.5
R16 Y.n1 Y.t2 36.818
R17 Y Y.n2 26.176
R18 Y.n0 Y.t1 14.021
R19 VGND.n0 VGND.t0 89.912
R20 VGND.n0 VGND.t1 78.487
R21 VGND VGND.n0 0.002
R22 B1.n0 B1.t0 510.919
R23 B1.n0 B1.t1 200.832
R24 B1 B1.n0 66.219
C0 Y B1 0.19fF
C1 A1 VPWR 0.07fF
C2 A1 a_116_351# 0.11fF
C3 VPWR a_227_47# 0.00fF
C4 a_227_47# a_116_351# 0.01fF
C5 A1 A2 0.07fF
C6 A2 a_227_47# 0.01fF
C7 Y A1 0.01fF
C8 Y a_227_47# 0.01fF
C9 VPWR a_116_351# 0.62fF
C10 VPWR A2 0.04fF
C11 A2 a_116_351# 0.09fF
C12 VPWR B1 0.03fF
C13 B1 a_116_351# 0.01fF
C14 A2 B1 0.03fF
C15 Y VPWR 0.10fF
C16 Y a_116_351# 0.15fF
C17 Y A2 0.06fF
.ends

