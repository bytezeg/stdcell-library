magic
tech sky130A
magscale 1 2
timestamp 1678771731
<< nwell >>
rect -38 315 498 998
<< nmos >>
rect 200 47 230 223
rect 312 47 342 223
<< pmos >>
rect 200 351 230 913
rect 312 351 342 913
<< ndiff >>
rect 118 170 200 223
rect 118 136 138 170
rect 172 136 200 170
rect 118 102 200 136
rect 118 68 138 102
rect 172 68 200 102
rect 118 47 200 68
rect 230 47 312 223
rect 342 170 424 223
rect 342 136 366 170
rect 400 136 424 170
rect 342 102 424 136
rect 342 68 366 102
rect 400 68 424 102
rect 342 47 424 68
<< pdiff >>
rect 110 892 200 913
rect 110 858 147 892
rect 181 858 200 892
rect 110 824 200 858
rect 110 790 147 824
rect 181 790 200 824
rect 110 756 200 790
rect 110 722 147 756
rect 181 722 200 756
rect 110 688 200 722
rect 110 654 147 688
rect 181 654 200 688
rect 110 620 200 654
rect 110 586 147 620
rect 181 586 200 620
rect 110 552 200 586
rect 110 518 147 552
rect 181 518 200 552
rect 110 484 200 518
rect 110 450 147 484
rect 181 450 200 484
rect 110 351 200 450
rect 230 892 312 913
rect 230 858 255 892
rect 289 858 312 892
rect 230 824 312 858
rect 230 790 255 824
rect 289 790 312 824
rect 230 756 312 790
rect 230 722 255 756
rect 289 722 312 756
rect 230 688 312 722
rect 230 654 255 688
rect 289 654 312 688
rect 230 620 312 654
rect 230 586 255 620
rect 289 586 312 620
rect 230 552 312 586
rect 230 518 255 552
rect 289 518 312 552
rect 230 484 312 518
rect 230 450 255 484
rect 289 450 312 484
rect 230 351 312 450
rect 342 892 424 913
rect 342 858 366 892
rect 400 858 424 892
rect 342 824 424 858
rect 342 790 366 824
rect 400 790 424 824
rect 342 756 424 790
rect 342 722 366 756
rect 400 722 424 756
rect 342 688 424 722
rect 342 654 366 688
rect 400 654 424 688
rect 342 620 424 654
rect 342 586 366 620
rect 400 586 424 620
rect 342 552 424 586
rect 342 518 366 552
rect 400 518 424 552
rect 342 484 424 518
rect 342 450 366 484
rect 400 450 424 484
rect 342 351 424 450
<< ndiffc >>
rect 138 136 172 170
rect 138 68 172 102
rect 366 136 400 170
rect 366 68 400 102
<< pdiffc >>
rect 147 858 181 892
rect 147 790 181 824
rect 147 722 181 756
rect 147 654 181 688
rect 147 586 181 620
rect 147 518 181 552
rect 147 450 181 484
rect 255 858 289 892
rect 255 790 289 824
rect 255 722 289 756
rect 255 654 289 688
rect 255 586 289 620
rect 255 518 289 552
rect 255 450 289 484
rect 366 858 400 892
rect 366 790 400 824
rect 366 722 400 756
rect 366 654 400 688
rect 366 586 400 620
rect 366 518 400 552
rect 366 450 400 484
<< psubdiff >>
rect 36 173 118 223
rect 36 139 56 173
rect 90 139 118 173
rect 36 105 118 139
rect 36 71 56 105
rect 90 71 118 105
rect 36 47 118 71
<< nsubdiff >>
rect 36 889 110 913
rect 36 855 52 889
rect 86 855 110 889
rect 36 821 110 855
rect 36 787 52 821
rect 86 787 110 821
rect 36 753 110 787
rect 36 719 52 753
rect 86 719 110 753
rect 36 685 110 719
rect 36 651 52 685
rect 86 651 110 685
rect 36 617 110 651
rect 36 583 52 617
rect 86 583 110 617
rect 36 549 110 583
rect 36 515 52 549
rect 86 515 110 549
rect 36 481 110 515
rect 36 447 52 481
rect 86 447 110 481
rect 36 351 110 447
<< psubdiffcont >>
rect 56 139 90 173
rect 56 71 90 105
<< nsubdiffcont >>
rect 52 855 86 889
rect 52 787 86 821
rect 52 719 86 753
rect 52 651 86 685
rect 52 583 86 617
rect 52 515 86 549
rect 52 447 86 481
<< poly >>
rect 200 913 230 939
rect 312 913 342 939
rect 200 314 230 351
rect 312 314 342 351
rect 80 304 230 314
rect 80 270 109 304
rect 143 270 177 304
rect 211 270 230 304
rect 80 260 230 270
rect 296 304 431 314
rect 296 270 313 304
rect 347 270 381 304
rect 415 270 431 304
rect 296 260 431 270
rect 200 223 230 260
rect 312 223 342 260
rect 200 21 230 47
rect 312 21 342 47
<< polycont >>
rect 109 270 143 304
rect 177 270 211 304
rect 313 270 347 304
rect 381 270 415 304
<< locali >>
rect 0 943 29 977
rect 63 943 121 977
rect 155 943 213 977
rect 247 943 305 977
rect 339 943 397 977
rect 431 943 460 977
rect 36 892 202 943
rect 36 889 147 892
rect 36 855 52 889
rect 86 858 147 889
rect 181 858 202 892
rect 86 855 202 858
rect 36 824 202 855
rect 36 821 147 824
rect 36 787 52 821
rect 86 790 147 821
rect 181 790 202 824
rect 86 787 202 790
rect 36 756 202 787
rect 36 753 147 756
rect 36 719 52 753
rect 86 722 147 753
rect 181 722 202 756
rect 86 719 202 722
rect 36 688 202 719
rect 36 685 147 688
rect 36 651 52 685
rect 86 654 147 685
rect 181 654 202 688
rect 86 651 202 654
rect 36 620 202 651
rect 36 617 147 620
rect 36 583 52 617
rect 86 586 147 617
rect 181 586 202 620
rect 86 583 202 586
rect 36 552 202 583
rect 36 549 147 552
rect 36 515 52 549
rect 86 518 147 549
rect 181 518 202 552
rect 86 515 202 518
rect 36 484 202 515
rect 36 481 147 484
rect 36 447 52 481
rect 86 450 147 481
rect 181 450 202 484
rect 86 447 202 450
rect 36 440 202 447
rect 245 892 294 908
rect 245 858 255 892
rect 289 858 294 892
rect 245 824 294 858
rect 245 790 255 824
rect 289 790 294 824
rect 245 756 294 790
rect 245 722 255 756
rect 289 722 294 756
rect 245 688 294 722
rect 245 654 255 688
rect 289 654 294 688
rect 245 620 294 654
rect 245 586 255 620
rect 289 586 294 620
rect 245 552 294 586
rect 245 518 255 552
rect 289 518 294 552
rect 245 484 294 518
rect 245 450 255 484
rect 289 450 294 484
rect 245 434 294 450
rect 366 892 400 943
rect 366 824 400 858
rect 366 756 400 790
rect 366 688 400 722
rect 366 620 400 654
rect 366 552 400 586
rect 366 484 400 518
rect 366 434 400 450
rect 109 304 211 387
rect 143 270 177 304
rect 109 254 211 270
rect 245 186 279 434
rect 313 304 415 388
rect 347 270 381 304
rect 313 254 415 270
rect 36 173 172 186
rect 36 139 56 173
rect 90 170 172 173
rect 90 139 138 170
rect 36 136 138 139
rect 245 170 400 186
rect 245 148 366 170
rect 36 105 172 136
rect 36 71 56 105
rect 90 102 172 105
rect 90 71 138 102
rect 36 68 138 71
rect 36 17 172 68
rect 365 136 366 148
rect 365 102 400 136
rect 365 68 366 102
rect 365 51 400 68
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 943 63 977
rect 121 943 155 977
rect 213 943 247 977
rect 305 943 339 977
rect 397 943 431 977
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 977 460 1000
rect 0 943 29 977
rect 63 943 121 977
rect 155 943 213 977
rect 247 943 305 977
rect 339 943 397 977
rect 431 943 460 977
rect 0 920 460 943
rect 0 17 460 40
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -40 460 -17
<< labels >>
flabel metal1 s 221 943 255 977 0 FreeSans 240 0 0 0 VPWR
port 3 nsew power bidirectional
flabel metal1 s 221 -17 255 17 0 FreeSans 240 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 121 343 155 377 0 FreeSans 240 0 0 0 A1
port 0 nsew signal input
flabel locali s 351 343 385 377 0 FreeSans 240 0 0 0 B1
port 1 nsew signal input
flabel locali s 245 343 279 377 0 FreeSans 240 0 0 0 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 460 960
string LEFclass CORE
string LEForigin 0 0
<< end >>
