magic
tech sky130A
magscale 1 2
timestamp 1682099520
<< nwell >>
rect -38 316 866 998
rect 0 315 866 316
<< nmos >>
rect 195 47 225 223
rect 349 47 379 223
rect 503 47 533 223
rect 657 47 687 223
<< pmos >>
rect 195 351 225 913
rect 349 351 379 913
rect 503 351 533 913
rect 657 351 687 913
<< ndiff >>
rect 115 173 195 223
rect 115 139 138 173
rect 172 139 195 173
rect 115 105 195 139
rect 115 71 138 105
rect 172 71 195 105
rect 115 47 195 71
rect 225 105 349 223
rect 225 71 236 105
rect 270 71 304 105
rect 338 71 349 105
rect 225 47 349 71
rect 379 173 503 223
rect 379 139 422 173
rect 456 139 503 173
rect 379 105 503 139
rect 379 71 422 105
rect 456 71 503 105
rect 379 47 503 71
rect 533 47 657 223
rect 687 173 767 223
rect 687 139 710 173
rect 744 139 767 173
rect 687 105 767 139
rect 687 71 710 105
rect 744 71 767 105
rect 687 47 767 71
<< pdiff >>
rect 115 889 195 913
rect 115 855 138 889
rect 172 855 195 889
rect 115 821 195 855
rect 115 787 138 821
rect 172 787 195 821
rect 115 753 195 787
rect 115 719 138 753
rect 172 719 195 753
rect 115 685 195 719
rect 115 651 138 685
rect 172 651 195 685
rect 115 617 195 651
rect 115 583 138 617
rect 172 583 195 617
rect 115 549 195 583
rect 115 515 138 549
rect 172 515 195 549
rect 115 481 195 515
rect 115 447 138 481
rect 172 447 195 481
rect 115 351 195 447
rect 225 351 349 913
rect 379 889 503 913
rect 379 855 423 889
rect 457 855 503 889
rect 379 821 503 855
rect 379 787 423 821
rect 457 787 503 821
rect 379 753 503 787
rect 379 719 423 753
rect 457 719 503 753
rect 379 685 503 719
rect 379 651 423 685
rect 457 651 503 685
rect 379 617 503 651
rect 379 583 423 617
rect 457 583 503 617
rect 379 549 503 583
rect 379 515 423 549
rect 457 515 503 549
rect 379 481 503 515
rect 379 447 423 481
rect 457 447 503 481
rect 379 351 503 447
rect 533 889 657 913
rect 533 855 544 889
rect 578 855 612 889
rect 646 855 657 889
rect 533 821 657 855
rect 533 787 544 821
rect 578 787 612 821
rect 646 787 657 821
rect 533 753 657 787
rect 533 719 544 753
rect 578 719 612 753
rect 646 719 657 753
rect 533 685 657 719
rect 533 651 544 685
rect 578 651 612 685
rect 646 651 657 685
rect 533 617 657 651
rect 533 583 544 617
rect 578 583 612 617
rect 646 583 657 617
rect 533 351 657 583
rect 687 889 767 913
rect 687 855 710 889
rect 744 855 767 889
rect 687 821 767 855
rect 687 787 710 821
rect 744 787 767 821
rect 687 753 767 787
rect 687 719 710 753
rect 744 719 767 753
rect 687 685 767 719
rect 687 651 710 685
rect 744 651 767 685
rect 687 617 767 651
rect 687 583 710 617
rect 744 583 767 617
rect 687 549 767 583
rect 687 515 710 549
rect 744 515 767 549
rect 687 481 767 515
rect 687 447 710 481
rect 744 447 767 481
rect 687 351 767 447
<< ndiffc >>
rect 138 139 172 173
rect 138 71 172 105
rect 236 71 270 105
rect 304 71 338 105
rect 422 139 456 173
rect 422 71 456 105
rect 710 139 744 173
rect 710 71 744 105
<< pdiffc >>
rect 138 855 172 889
rect 138 787 172 821
rect 138 719 172 753
rect 138 651 172 685
rect 138 583 172 617
rect 138 515 172 549
rect 138 447 172 481
rect 423 855 457 889
rect 423 787 457 821
rect 423 719 457 753
rect 423 651 457 685
rect 423 583 457 617
rect 423 515 457 549
rect 423 447 457 481
rect 544 855 578 889
rect 612 855 646 889
rect 544 787 578 821
rect 612 787 646 821
rect 544 719 578 753
rect 612 719 646 753
rect 544 651 578 685
rect 612 651 646 685
rect 544 583 578 617
rect 612 583 646 617
rect 710 855 744 889
rect 710 787 744 821
rect 710 719 744 753
rect 710 651 744 685
rect 710 583 744 617
rect 710 515 744 549
rect 710 447 744 481
<< psubdiff >>
rect 36 173 115 223
rect 36 139 59 173
rect 93 139 115 173
rect 36 105 115 139
rect 36 71 59 105
rect 93 71 115 105
rect 36 47 115 71
<< nsubdiff >>
rect 36 889 115 913
rect 36 855 59 889
rect 93 855 115 889
rect 36 821 115 855
rect 36 787 59 821
rect 93 787 115 821
rect 36 753 115 787
rect 36 719 59 753
rect 93 719 115 753
rect 36 685 115 719
rect 36 651 59 685
rect 93 651 115 685
rect 36 617 115 651
rect 36 583 59 617
rect 93 583 115 617
rect 36 549 115 583
rect 36 515 59 549
rect 93 515 115 549
rect 36 481 115 515
rect 36 447 59 481
rect 93 447 115 481
rect 36 351 115 447
<< psubdiffcont >>
rect 59 139 93 173
rect 59 71 93 105
<< nsubdiffcont >>
rect 59 855 93 889
rect 59 787 93 821
rect 59 719 93 753
rect 59 651 93 685
rect 59 583 93 617
rect 59 515 93 549
rect 59 447 93 481
<< poly >>
rect 195 913 225 939
rect 349 913 379 939
rect 503 913 533 939
rect 657 913 687 939
rect 195 314 225 351
rect 349 314 379 351
rect 503 314 533 351
rect 657 314 687 351
rect 61 304 225 314
rect 61 270 77 304
rect 111 270 145 304
rect 179 270 225 304
rect 61 260 225 270
rect 267 304 401 314
rect 267 270 283 304
rect 317 270 351 304
rect 385 270 401 304
rect 267 260 401 270
rect 443 304 579 314
rect 443 270 459 304
rect 493 270 527 304
rect 561 270 579 304
rect 443 260 579 270
rect 657 304 791 314
rect 657 270 673 304
rect 707 270 741 304
rect 775 270 791 304
rect 657 260 791 270
rect 195 223 225 260
rect 349 223 379 260
rect 503 223 533 260
rect 657 223 687 260
rect 195 21 225 47
rect 349 21 379 47
rect 503 21 533 47
rect 657 21 687 47
<< polycont >>
rect 77 270 111 304
rect 145 270 179 304
rect 283 270 317 304
rect 351 270 385 304
rect 459 270 493 304
rect 527 270 561 304
rect 673 270 707 304
rect 741 270 775 304
<< locali >>
rect 0 943 29 977
rect 63 943 121 977
rect 155 943 213 977
rect 247 943 305 977
rect 339 943 397 977
rect 431 943 489 977
rect 523 943 581 977
rect 615 943 673 977
rect 707 943 765 977
rect 799 943 828 977
rect 59 889 172 943
rect 93 855 138 889
rect 59 821 172 855
rect 93 787 138 821
rect 59 753 172 787
rect 93 719 138 753
rect 59 685 172 719
rect 93 651 138 685
rect 59 617 172 651
rect 93 583 138 617
rect 59 549 172 583
rect 93 515 138 549
rect 59 481 172 515
rect 93 447 138 481
rect 59 431 172 447
rect 423 889 457 909
rect 423 821 457 855
rect 423 753 457 787
rect 423 685 457 719
rect 423 617 457 651
rect 423 549 457 583
rect 544 889 646 943
rect 578 855 612 889
rect 544 821 646 855
rect 578 787 612 821
rect 544 753 646 787
rect 578 719 612 753
rect 544 685 646 719
rect 578 651 612 685
rect 544 617 646 651
rect 578 583 612 617
rect 544 567 646 583
rect 710 889 744 909
rect 710 821 744 855
rect 710 753 744 787
rect 710 685 744 719
rect 710 617 744 651
rect 423 481 457 515
rect 710 549 744 583
rect 710 481 744 515
rect 457 447 710 481
rect 423 431 744 447
rect 77 304 179 386
rect 111 270 145 304
rect 77 254 179 270
rect 283 304 385 386
rect 317 270 351 304
rect 283 254 385 270
rect 459 304 561 386
rect 493 270 527 304
rect 459 254 561 270
rect 595 201 629 431
rect 673 304 781 386
rect 707 270 741 304
rect 775 270 781 304
rect 673 254 781 270
rect 59 173 93 190
rect 59 105 93 139
rect 59 17 93 71
rect 138 173 456 190
rect 172 156 422 173
rect 138 105 172 139
rect 595 173 744 201
rect 595 167 710 173
rect 422 105 456 139
rect 138 51 172 71
rect 220 71 236 105
rect 270 71 304 105
rect 338 71 354 105
rect 220 17 354 71
rect 422 51 456 71
rect 710 105 744 139
rect 710 51 744 71
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 943 63 977
rect 121 943 155 977
rect 213 943 247 977
rect 305 943 339 977
rect 397 943 431 977
rect 489 943 523 977
rect 581 943 615 977
rect 673 943 707 977
rect 765 943 799 977
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 977 828 1000
rect 0 943 29 977
rect 63 943 121 977
rect 155 943 213 977
rect 247 943 305 977
rect 339 943 397 977
rect 431 943 489 977
rect 523 943 581 977
rect 615 943 673 977
rect 707 943 765 977
rect 799 943 828 977
rect 0 920 828 943
rect 0 17 828 40
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -40 828 -17
<< labels >>
flabel locali s 305 343 339 377 0 FreeSans 240 0 0 0 A1
port 1 nsew signal input
flabel locali s 489 343 523 377 0 FreeSans 240 0 0 0 B1
port 2 nsew
flabel locali s 595 263 629 297 0 FreeSans 240 0 0 0 Y
port 4 nsew signal output
flabel metal1 s 397 943 431 977 0 FreeSans 240 0 0 0 VPWR
port 5 nsew power bidirectional
flabel locali s 716 343 750 377 0 FreeSans 240 0 0 0 C1
port 3 nsew signal input
flabel locali s 121 343 155 377 0 FreeSans 240 0 0 0 A2
port 0 nsew signal input
flabel metal1 s 397 -17 431 17 0 FreeSans 240 0 0 0 VGND
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 828 960
string LEFclass CORE
string LEForigin 0 0
<< end >>
