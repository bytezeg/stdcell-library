magic
tech sky130A
magscale 1 2
timestamp 1678775228
<< nwell >>
rect -38 314 406 998
<< nmos >>
rect 213 47 243 223
<< pmos >>
rect 213 351 243 913
<< ndiff >>
rect 125 157 213 223
rect 125 123 152 157
rect 186 123 213 157
rect 125 89 213 123
rect 125 55 152 89
rect 186 55 213 89
rect 125 47 213 55
rect 243 157 332 223
rect 243 123 268 157
rect 302 123 332 157
rect 243 89 332 123
rect 243 55 268 89
rect 302 55 332 89
rect 243 47 332 55
<< pdiff >>
rect 125 905 213 913
rect 125 871 152 905
rect 186 871 213 905
rect 125 837 213 871
rect 125 803 152 837
rect 186 803 213 837
rect 125 769 213 803
rect 125 735 152 769
rect 186 735 213 769
rect 125 701 213 735
rect 125 667 152 701
rect 186 667 213 701
rect 125 633 213 667
rect 125 599 152 633
rect 186 599 213 633
rect 125 565 213 599
rect 125 531 152 565
rect 186 531 213 565
rect 125 351 213 531
rect 243 905 332 913
rect 243 871 269 905
rect 304 871 332 905
rect 243 837 332 871
rect 243 803 268 837
rect 304 803 332 837
rect 243 769 332 803
rect 243 735 268 769
rect 304 735 332 769
rect 243 701 332 735
rect 243 667 268 701
rect 304 667 332 701
rect 243 633 332 667
rect 243 599 268 633
rect 304 599 332 633
rect 243 565 332 599
rect 243 531 268 565
rect 304 531 332 565
rect 243 351 332 531
<< ndiffc >>
rect 152 123 186 157
rect 152 55 186 89
rect 268 123 302 157
rect 268 55 302 89
<< pdiffc >>
rect 152 871 186 905
rect 152 803 186 837
rect 152 735 186 769
rect 152 667 186 701
rect 152 599 186 633
rect 152 531 186 565
rect 269 871 304 905
rect 268 803 304 837
rect 268 735 304 769
rect 268 667 304 701
rect 268 599 304 633
rect 268 531 304 565
<< psubdiff >>
rect 36 157 125 223
rect 36 123 63 157
rect 97 123 125 157
rect 36 89 125 123
rect 36 55 63 89
rect 97 55 125 89
rect 36 47 125 55
<< nsubdiff >>
rect 36 905 125 913
rect 36 871 63 905
rect 97 871 125 905
rect 36 837 125 871
rect 36 803 63 837
rect 97 803 125 837
rect 36 769 125 803
rect 36 735 63 769
rect 97 735 125 769
rect 36 701 125 735
rect 36 667 63 701
rect 97 667 125 701
rect 36 633 125 667
rect 36 599 63 633
rect 97 599 125 633
rect 36 565 125 599
rect 36 531 63 565
rect 97 531 125 565
rect 36 351 125 531
<< psubdiffcont >>
rect 63 123 97 157
rect 63 55 97 89
<< nsubdiffcont >>
rect 63 871 97 905
rect 63 803 97 837
rect 63 735 97 769
rect 63 667 97 701
rect 63 599 97 633
rect 63 531 97 565
<< poly >>
rect 213 913 243 939
rect 213 314 243 351
rect 79 304 243 314
rect 79 270 95 304
rect 129 270 163 304
rect 197 270 243 304
rect 79 260 243 270
rect 213 223 243 260
rect 213 21 243 47
<< polycont >>
rect 95 270 129 304
rect 163 270 197 304
<< locali >>
rect 0 943 29 977
rect 63 943 121 977
rect 155 943 213 977
rect 247 943 305 977
rect 339 943 368 977
rect 63 905 202 943
rect 97 871 152 905
rect 63 837 186 871
rect 97 803 152 837
rect 63 769 186 803
rect 97 735 152 769
rect 63 701 186 735
rect 97 667 152 701
rect 63 633 186 667
rect 97 599 152 633
rect 63 565 186 599
rect 97 531 152 565
rect 63 502 186 531
rect 252 871 269 905
rect 304 871 320 905
rect 252 837 320 871
rect 252 803 268 837
rect 304 803 320 837
rect 252 769 320 803
rect 252 735 268 769
rect 304 735 320 769
rect 252 701 320 735
rect 252 667 268 701
rect 304 667 320 701
rect 252 633 320 667
rect 252 599 268 633
rect 304 599 320 633
rect 252 565 320 599
rect 252 531 268 565
rect 304 531 320 565
rect 78 304 213 460
rect 78 270 95 304
rect 129 270 163 304
rect 197 270 213 304
rect 78 220 213 270
rect 63 157 202 173
rect 97 123 152 157
rect 186 123 202 157
rect 63 89 202 123
rect 97 55 152 89
rect 186 55 202 89
rect 63 17 202 55
rect 252 157 320 531
rect 252 123 268 157
rect 302 123 320 157
rect 252 89 320 123
rect 252 55 268 89
rect 302 55 320 89
rect 252 52 320 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< viali >>
rect 29 943 63 977
rect 121 943 155 977
rect 213 943 247 977
rect 305 943 339 977
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 977 368 1000
rect 0 943 29 977
rect 63 943 121 977
rect 155 943 213 977
rect 247 943 305 977
rect 339 943 368 977
rect 0 920 368 943
rect 0 17 368 40
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -40 368 -17
<< labels >>
flabel metal1 s 0 920 368 1000 0 FreeSans 240 0 0 0 VPWR
port 2 nsew power bidirectional
flabel metal1 s 0 -40 368 40 0 FreeSans 240 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 121 343 155 377 0 FreeSans 240 0 0 0 A
port 0 nsew signal input
flabel locali s 254 343 288 377 0 FreeSans 240 0 0 0 Y
port 1 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 368 960
string LEFclass CORE
string LEForigin 0 0
<< end >>
