magic
tech sky130A
magscale 1 2
timestamp 1678760939
<< nwell >>
rect -38 315 858 998
<< nmos >>
rect 195 47 225 223
rect 349 47 379 223
rect 503 47 533 223
rect 657 47 687 223
<< pmos >>
rect 195 351 225 913
rect 349 351 379 913
rect 503 351 533 913
rect 657 351 687 913
<< ndiff >>
rect 115 173 195 223
rect 115 139 138 173
rect 172 139 195 173
rect 115 105 195 139
rect 115 71 138 105
rect 172 71 195 105
rect 115 47 195 71
rect 225 47 349 223
rect 379 173 503 223
rect 379 139 424 173
rect 458 139 503 173
rect 379 105 503 139
rect 379 71 424 105
rect 458 71 503 105
rect 379 47 503 71
rect 533 47 657 223
rect 687 169 767 223
rect 687 135 710 169
rect 744 135 767 169
rect 687 101 767 135
rect 687 67 710 101
rect 744 67 767 101
rect 687 47 767 67
<< pdiff >>
rect 115 821 195 913
rect 115 787 138 821
rect 172 787 195 821
rect 115 753 195 787
rect 115 719 138 753
rect 172 719 195 753
rect 115 685 195 719
rect 115 651 138 685
rect 172 651 195 685
rect 115 617 195 651
rect 115 583 138 617
rect 172 583 195 617
rect 115 549 195 583
rect 115 515 138 549
rect 172 515 195 549
rect 115 351 195 515
rect 225 821 349 913
rect 225 787 270 821
rect 304 787 349 821
rect 225 753 349 787
rect 225 719 270 753
rect 304 719 349 753
rect 225 685 349 719
rect 225 651 270 685
rect 304 651 349 685
rect 225 617 349 651
rect 225 583 270 617
rect 304 583 349 617
rect 225 549 349 583
rect 225 515 270 549
rect 304 515 349 549
rect 225 351 349 515
rect 379 821 503 913
rect 379 787 418 821
rect 452 787 503 821
rect 379 753 503 787
rect 379 719 418 753
rect 452 719 503 753
rect 379 685 503 719
rect 379 651 418 685
rect 452 651 503 685
rect 379 617 503 651
rect 379 583 418 617
rect 452 583 503 617
rect 379 549 503 583
rect 379 515 418 549
rect 452 515 503 549
rect 379 351 503 515
rect 533 821 657 913
rect 533 787 578 821
rect 612 787 657 821
rect 533 753 657 787
rect 533 719 578 753
rect 612 719 657 753
rect 533 685 657 719
rect 533 651 578 685
rect 612 651 657 685
rect 533 617 657 651
rect 533 583 578 617
rect 612 583 657 617
rect 533 549 657 583
rect 533 515 578 549
rect 612 515 657 549
rect 533 351 657 515
rect 687 821 775 913
rect 687 787 698 821
rect 732 787 775 821
rect 687 753 775 787
rect 687 719 698 753
rect 732 719 775 753
rect 687 685 775 719
rect 687 651 698 685
rect 732 651 775 685
rect 687 617 775 651
rect 687 583 698 617
rect 732 583 775 617
rect 687 549 775 583
rect 687 515 698 549
rect 732 515 775 549
rect 687 481 775 515
rect 687 447 698 481
rect 732 447 775 481
rect 687 351 775 447
<< ndiffc >>
rect 138 139 172 173
rect 138 71 172 105
rect 424 139 458 173
rect 424 71 458 105
rect 710 135 744 169
rect 710 67 744 101
<< pdiffc >>
rect 138 787 172 821
rect 138 719 172 753
rect 138 651 172 685
rect 138 583 172 617
rect 138 515 172 549
rect 270 787 304 821
rect 270 719 304 753
rect 270 651 304 685
rect 270 583 304 617
rect 270 515 304 549
rect 418 787 452 821
rect 418 719 452 753
rect 418 651 452 685
rect 418 583 452 617
rect 418 515 452 549
rect 578 787 612 821
rect 578 719 612 753
rect 578 651 612 685
rect 578 583 612 617
rect 578 515 612 549
rect 698 787 732 821
rect 698 719 732 753
rect 698 651 732 685
rect 698 583 732 617
rect 698 515 732 549
rect 698 447 732 481
<< psubdiff >>
rect 36 173 115 223
rect 36 139 59 173
rect 93 139 115 173
rect 36 105 115 139
rect 36 71 59 105
rect 93 71 115 105
rect 36 47 115 71
<< nsubdiff >>
rect 36 821 115 913
rect 36 787 59 821
rect 93 787 115 821
rect 36 753 115 787
rect 36 719 59 753
rect 93 719 115 753
rect 36 685 115 719
rect 36 651 59 685
rect 93 651 115 685
rect 36 617 115 651
rect 36 583 59 617
rect 93 583 115 617
rect 36 549 115 583
rect 36 515 59 549
rect 93 515 115 549
rect 36 351 115 515
<< psubdiffcont >>
rect 59 139 93 173
rect 59 71 93 105
<< nsubdiffcont >>
rect 59 787 93 821
rect 59 719 93 753
rect 59 651 93 685
rect 59 583 93 617
rect 59 515 93 549
<< poly >>
rect 195 913 225 939
rect 349 913 379 939
rect 503 913 533 939
rect 657 913 687 939
rect 195 314 225 351
rect 349 314 379 351
rect 503 314 533 351
rect 657 314 687 351
rect 61 304 225 314
rect 61 270 77 304
rect 111 270 145 304
rect 179 270 225 304
rect 61 260 225 270
rect 267 304 401 314
rect 267 270 283 304
rect 317 270 351 304
rect 385 270 401 304
rect 267 260 401 270
rect 443 304 579 314
rect 443 270 459 304
rect 493 270 527 304
rect 561 270 579 304
rect 443 260 579 270
rect 657 304 797 314
rect 657 270 679 304
rect 713 270 747 304
rect 781 270 797 304
rect 657 260 797 270
rect 195 223 225 260
rect 349 223 379 260
rect 503 223 533 260
rect 657 223 687 260
rect 195 21 225 47
rect 349 21 379 47
rect 503 21 533 47
rect 657 21 687 47
<< polycont >>
rect 77 270 111 304
rect 145 270 179 304
rect 283 270 317 304
rect 351 270 385 304
rect 459 270 493 304
rect 527 270 561 304
rect 679 270 713 304
rect 747 270 781 304
<< locali >>
rect 0 943 29 977
rect 63 943 121 977
rect 155 943 213 977
rect 247 943 305 977
rect 339 943 397 977
rect 431 943 489 977
rect 523 943 581 977
rect 615 943 673 977
rect 707 943 765 977
rect 799 943 828 977
rect 59 821 93 943
rect 59 753 93 787
rect 59 685 93 719
rect 59 617 93 651
rect 59 549 93 583
rect 59 494 93 515
rect 138 821 172 905
rect 138 753 172 787
rect 138 685 172 719
rect 138 617 172 651
rect 138 549 172 583
rect 138 465 172 515
rect 270 821 304 943
rect 270 753 304 787
rect 270 685 304 719
rect 270 617 304 651
rect 270 549 304 583
rect 270 499 304 515
rect 418 871 732 905
rect 418 821 452 871
rect 418 753 452 787
rect 418 685 452 719
rect 418 617 452 651
rect 418 549 452 583
rect 418 465 452 515
rect 578 821 629 837
rect 612 787 629 821
rect 578 753 629 787
rect 612 719 629 753
rect 578 685 629 719
rect 612 651 629 685
rect 578 617 629 651
rect 612 583 629 617
rect 578 549 629 583
rect 612 515 629 549
rect 578 499 629 515
rect 138 431 452 465
rect 77 304 179 382
rect 111 270 145 304
rect 77 254 179 270
rect 283 304 385 382
rect 317 270 351 304
rect 283 254 385 270
rect 459 304 561 382
rect 493 270 527 304
rect 459 254 561 270
rect 595 211 629 499
rect 698 821 732 871
rect 698 753 732 787
rect 698 685 732 719
rect 698 617 732 651
rect 698 549 732 583
rect 698 481 732 515
rect 698 431 732 447
rect 679 304 781 382
rect 713 270 747 304
rect 679 254 781 270
rect 41 173 184 189
rect 41 139 59 173
rect 93 139 138 173
rect 172 139 184 173
rect 41 105 184 139
rect 41 71 59 105
rect 93 71 138 105
rect 172 71 184 105
rect 41 17 184 71
rect 424 177 629 211
rect 424 173 458 177
rect 424 105 458 139
rect 424 55 458 71
rect 710 169 744 185
rect 710 101 744 135
rect 710 17 744 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 943 63 977
rect 121 943 155 977
rect 213 943 247 977
rect 305 943 339 977
rect 397 943 431 977
rect 489 943 523 977
rect 581 943 615 977
rect 673 943 707 977
rect 765 943 799 977
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 977 828 1000
rect 0 943 29 977
rect 63 943 121 977
rect 155 943 213 977
rect 247 943 305 977
rect 339 943 397 977
rect 431 943 489 977
rect 523 943 581 977
rect 615 943 673 977
rect 707 943 765 977
rect 799 943 828 977
rect 0 920 828 943
rect 0 17 828 40
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -40 828 -17
<< labels >>
flabel locali s 121 343 155 377 0 FreeSans 240 0 0 0 A2
port 0 nsew signal input
flabel locali s 305 343 339 377 0 FreeSans 240 0 0 0 A1
port 1 nsew signal input
flabel locali s 489 343 523 377 0 FreeSans 240 0 0 0 B1
port 2 nsew signal input
flabel locali s 714 343 748 377 0 FreeSans 240 0 0 0 B2
port 3 nsew signal input
flabel locali s 595 280 629 314 0 FreeSans 240 0 0 0 Y
port 4 nsew signal output
flabel metal1 s 339 943 397 977 0 FreeSans 240 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 431 -17 489 17 0 FreeSans 240 0 0 0 VGND
port 6 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 828 960
string LEFclass CORE
string LEForigin 0 0
<< end >>
