* NGSPICE file created from thesis_buff.ext - technology: sky130A

.subckt thesis_buff A1 Y VPWR VGND
X0 Y.t1 a_110_351# VGND.t1 VGND sky130_fd_pr__nfet_01v8 ad=0.3608 pd=2.58 as=0.1804 ps=1.29 w=0.88 l=0.15
X1 VGND.t0 A1.t0 a_110_351# VGND sky130_fd_pr__nfet_01v8 ad=0.1804 pd=1.29 as=0.3608 ps=2.58 w=0.88 l=0.15
X2 Y.t0 a_110_351# VPWR.t3 VPWR.t2 sky130_fd_pr__pfet_01v8 ad=1.1521 pd=6.44 as=0.57605 ps=3.22 w=2.81 l=0.15
X3 VPWR.t1 A1.t1 a_110_351# VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.57605 pd=3.22 as=1.2645 ps=6.52 w=2.81 l=0.15
R0 VGND VGND.n0 65.136
R1 VGND.n0 VGND.t1 27.954
R2 VGND.n0 VGND.t0 27.954
R3 Y Y.t0 151.337
R4 Y Y.t1 132.97
R5 A1.n0 A1.t1 510.919
R6 A1.n0 A1.t0 200.832
R7 A1 A1.n0 70.149
R8 VPWR.n2 VPWR.t0 271.474
R9 VPWR.t0 VPWR.t2 155.783
R10 VPWR.n1 VPWR.n0 93.649
R11 VPWR.n0 VPWR.t1 14.722
R12 VPWR.n0 VPWR.t3 14.021
R13 VPWR VPWR.n2 4.767
R14 VPWR VPWR.n1 0.33
C0 Y A1 0.00fF
C1 VPWR Y 0.18fF
C2 VPWR A1 0.06fF
C3 a_110_351# Y 0.17fF
C4 a_110_351# A1 0.32fF
C5 VPWR a_110_351# 0.46fF
.ends

