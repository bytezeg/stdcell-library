magic
tech sky130A
timestamp 1670805011
<< error_p >>
rect 80 65 95 66
rect 80 23 95 24
<< nwell >>
rect 0 112 145 347
<< nmos >>
rect 80 24 95 65
<< pmos >>
rect 80 130 95 315
<< ndiff >>
rect 47 53 80 65
rect 47 36 54 53
rect 71 36 80 53
rect 47 24 80 36
rect 95 53 125 65
rect 95 36 104 53
rect 121 36 125 53
rect 95 24 125 36
<< pdiff >>
rect 47 303 80 315
rect 47 286 54 303
rect 71 286 80 303
rect 47 269 80 286
rect 47 252 54 269
rect 71 252 80 269
rect 47 235 80 252
rect 47 218 54 235
rect 71 218 80 235
rect 47 201 80 218
rect 47 184 54 201
rect 71 184 80 201
rect 47 167 80 184
rect 47 150 54 167
rect 71 150 80 167
rect 47 130 80 150
rect 95 303 127 315
rect 95 286 104 303
rect 121 286 127 303
rect 95 269 127 286
rect 95 252 104 269
rect 121 252 127 269
rect 95 235 127 252
rect 95 218 104 235
rect 121 218 127 235
rect 95 201 127 218
rect 95 184 104 201
rect 121 184 127 201
rect 95 167 127 184
rect 95 150 104 167
rect 121 150 127 167
rect 95 130 127 150
<< ndiffc >>
rect 54 36 71 53
rect 104 36 121 53
<< pdiffc >>
rect 54 286 71 303
rect 54 252 71 269
rect 54 218 71 235
rect 54 184 71 201
rect 54 150 71 167
rect 104 286 121 303
rect 104 252 121 269
rect 104 218 121 235
rect 104 184 121 201
rect 104 150 121 167
<< psubdiff >>
rect 8 53 47 65
rect 8 36 20 53
rect 37 36 47 53
rect 8 24 47 36
rect 17 -8 34 24
<< nsubdiff >>
rect 18 303 47 315
rect 18 286 20 303
rect 37 286 47 303
rect 18 269 47 286
rect 18 252 20 269
rect 37 252 47 269
rect 18 235 47 252
rect 18 218 20 235
rect 37 218 47 235
rect 18 201 47 218
rect 18 184 20 201
rect 37 184 47 201
rect 18 167 47 184
rect 18 150 20 167
rect 37 150 47 167
rect 18 130 47 150
<< psubdiffcont >>
rect 20 36 37 53
<< nsubdiffcont >>
rect 20 286 37 303
rect 20 252 37 269
rect 20 218 37 235
rect 20 184 37 201
rect 20 150 37 167
<< poly >>
rect 80 315 95 328
rect 80 111 95 130
rect 0 106 95 111
rect 0 89 8 106
rect 25 89 95 106
rect 0 84 95 89
rect 80 65 95 84
rect 80 11 95 24
<< polycont >>
rect 8 89 25 106
<< locali >>
rect 20 311 37 327
rect 12 303 79 311
rect 12 286 20 303
rect 37 286 54 303
rect 71 286 79 303
rect 12 269 79 286
rect 12 252 20 269
rect 37 252 54 269
rect 71 252 79 269
rect 12 235 79 252
rect 12 218 20 235
rect 37 218 54 235
rect 71 218 79 235
rect 12 201 79 218
rect 12 184 20 201
rect 37 184 54 201
rect 71 184 79 201
rect 12 167 79 184
rect 12 150 20 167
rect 37 150 54 167
rect 71 150 79 167
rect 12 130 79 150
rect 96 303 129 311
rect 96 286 104 303
rect 121 286 129 303
rect 96 269 129 286
rect 96 252 104 269
rect 121 252 129 269
rect 96 235 129 252
rect 96 218 104 235
rect 121 218 129 235
rect 96 201 129 218
rect 96 184 104 201
rect 121 184 129 201
rect 96 167 129 184
rect 96 150 104 167
rect 121 150 129 167
rect 96 106 129 150
rect 0 89 8 106
rect 25 89 33 106
rect 96 89 104 106
rect 121 89 129 106
rect 12 53 79 61
rect 12 36 20 53
rect 37 36 54 53
rect 71 36 79 53
rect 12 28 79 36
rect 96 53 129 89
rect 96 36 104 53
rect 121 36 129 53
rect 96 28 129 36
rect 17 9 34 28
<< viali >>
rect 20 327 37 344
rect 8 89 25 106
rect 104 89 121 106
rect 17 -8 34 9
<< metal1 >>
rect 0 344 145 347
rect 0 327 20 344
rect 37 327 145 344
rect 0 324 145 327
rect 0 273 145 287
rect 0 245 145 259
rect 0 217 145 231
rect 0 189 145 203
rect 0 161 145 175
rect 0 133 145 147
rect 0 106 145 119
rect 0 89 8 106
rect 25 105 104 106
rect 25 91 28 105
rect 101 91 104 105
rect 25 89 104 91
rect 121 105 145 106
rect 121 91 124 105
rect 121 89 145 91
rect 0 77 145 89
rect 0 49 145 63
rect 0 9 145 12
rect 0 -8 17 9
rect 34 -8 145 9
rect 0 -11 145 -8
<< end >>
