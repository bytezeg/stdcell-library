* NGSPICE file created from thesis_aoi22.ext - technology: sky130A

.subckt thesis_aoi22 A2 A1 B1 B2 Y VPWR VGND
X0 a_115_351# A1.t0 VPWR.t1 VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.8711 pd=3.43 as=0.8711 ps=3.43 w=2.81 l=0.15
X1 Y.t0 A1.t1 a_225_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2728 pd=1.5 as=0.2728 ps=1.5 w=0.88 l=0.15
X2 a_533_47# B1.t0 Y.t1 VGND sky130_fd_pr__nfet_01v8 ad=0.2728 pd=1.5 as=0.2728 ps=1.5 w=0.88 l=0.15
X3 Y.t2 B1.t1 a_115_351# VPWR.t2 sky130_fd_pr__pfet_01v8 ad=0.8711 pd=3.43 as=0.8711 ps=3.43 w=2.81 l=0.15
X4 a_115_351# B2.t0 Y.t3 VPWR.t3 sky130_fd_pr__pfet_01v8 ad=1.2364 pd=6.5 as=0.8711 ps=3.43 w=2.81 l=0.15
X5 VGND.t1 B2.t1 a_533_47# VGND sky130_fd_pr__nfet_01v8 ad=0.352 pd=2.56 as=0.2728 ps=1.5 w=0.88 l=0.15
X6 VPWR.t5 A2.t0 a_115_351# VPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.8711 pd=3.43 as=1.124 ps=6.42 w=2.81 l=0.15
X7 a_225_47# A2.t1 VGND.t0 VGND sky130_fd_pr__nfet_01v8 ad=0.2728 pd=1.5 as=0.352 ps=2.56 w=0.88 l=0.15
R0 A1.n0 A1.t0 510.919
R1 A1.n0 A1.t1 200.832
R2 A1 A1.n0 52.276
R3 VPWR.n1 VPWR.t4 308.904
R4 VPWR.t2 VPWR.t3 214.202
R5 VPWR.t0 VPWR.t2 214.202
R6 VPWR.t4 VPWR.t0 214.202
R7 VPWR.n1 VPWR.n0 146.914
R8 VPWR.n0 VPWR.t1 21.733
R9 VPWR.n0 VPWR.t5 21.733
R10 VPWR VPWR.n1 0.162
R11 Y Y.n0 167.415
R12 Y Y.n1 150.13
R13 Y.n1 Y.t1 42.272
R14 Y.n1 Y.t0 42.272
R15 Y.n0 Y.t3 21.733
R16 Y.n0 Y.t2 21.733
R17 VGND.n0 VGND.t1 115.333
R18 VGND.n0 VGND.t0 85.415
R19 VGND.n0 VGND 0.001
R20 B1.n0 B1.t1 510.919
R21 B1.n0 B1.t0 200.832
R22 B1 B1.n0 54.758
R23 B2.n0 B2.t0 510.919
R24 B2.n0 B2.t1 200.832
R25 B2 B2.n0 71.646
R26 A2.n0 A2.t0 510.919
R27 A2.n0 A2.t1 200.832
R28 A2 A2.n0 93.713
C0 a_115_351# B2 0.11fF
C1 VPWR B2 0.02fF
C2 B1 Y 0.16fF
C3 a_115_351# A1 0.10fF
C4 VPWR A1 0.04fF
C5 a_115_351# A2 0.11fF
C6 a_115_351# Y 0.36fF
C7 VPWR A2 0.06fF
C8 VPWR Y 0.04fF
C9 a_533_47# Y 0.06fF
C10 a_115_351# B1 0.06fF
C11 A1 a_225_47# 0.02fF
C12 B1 VPWR 0.01fF
C13 B1 a_533_47# 0.00fF
C14 Y a_225_47# 0.01fF
C15 a_115_351# VPWR 0.91fF
C16 a_115_351# a_533_47# 0.00fF
C17 B2 Y 0.08fF
C18 a_533_47# VPWR 0.00fF
C19 A2 A1 0.07fF
C20 A1 Y 0.01fF
C21 B1 B2 0.03fF
C22 a_115_351# a_225_47# 0.02fF
C23 A2 Y 0.00fF
C24 B1 A1 0.07fF
C25 VPWR a_225_47# 0.00fF
.ends

