* NGSPICE file created from thesis_oai21.ext - technology: sky130A

.subckt thesis_oai21 A1 A2 B1 Y VPWR VGND
X0 Y.t2 A2.t0 a_216_351# VPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.765725 pd=3.355 as=0.765725 ps=3.355 w=2.81 l=0.15
X1 a_111_47# A2.t1 VGND.t1 VGND sky130_fd_pr__nfet_01v8 ad=0.2398 pd=1.425 as=0.2398 ps=1.425 w=0.88 l=0.15
X2 a_216_351# A1.t0 VPWR.t1 VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.765725 pd=3.355 as=1.05375 ps=6.37 w=2.81 l=0.15
X3 VPWR.t3 B1.t0 Y.t0 VPWR.t2 sky130_fd_pr__pfet_01v8 ad=1.05375 pd=6.37 as=0.765725 ps=3.355 w=2.81 l=0.15
X4 Y.t1 B1.t1 a_111_47# VGND sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.51 as=0.2398 ps=1.425 w=0.88 l=0.15
X5 VGND.t0 A1.t1 a_111_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2398 pd=1.425 as=0.33 ps=2.51 w=0.88 l=0.15
R0 A2.n0 A2.t0 510.919
R1 A2.n0 A2.t1 200.832
R2 A2 A2.n0 54.486
R3 Y Y.n0 243.65
R4 Y Y.t1 170.84
R5 Y.n0 Y.t0 19.279
R6 Y.n0 Y.t2 18.928
R7 VPWR.n4 VPWR.t1 376.553
R8 VPWR.n7 VPWR.n6 292.5
R9 VPWR.n9 VPWR.n8 292.5
R10 VPWR.t4 VPWR.t2 193.338
R11 VPWR.t0 VPWR.t4 193.338
R12 VPWR.n13 VPWR.t0 182.21
R13 VPWR.n0 VPWR.t3 134.107
R14 VPWR.n15 VPWR.n14 126.755
R15 VPWR.n7 VPWR.n5 92.5
R16 VPWR.n9 VPWR.n2 92.5
R17 VPWR.n11 VPWR.n10 92.5
R18 VPWR.n4 VPWR.n3 92.5
R19 VPWR.n2 VPWR.n1 34.255
R20 VPWR.n14 VPWR.n13 29.123
R21 VPWR.n16 VPWR.n15 11.426
R22 VPWR.n11 VPWR.n9 7.134
R23 VPWR.n9 VPWR.n7 7.134
R24 VPWR.n7 VPWR.n4 7.134
R25 VPWR.n15 VPWR.n12 4.361
R26 VPWR.n12 VPWR.n11 2.708
R27 VPWR VPWR.n16 0.61
R28 VPWR VPWR.n0 0.079
R29 VGND VGND.n0 67.584
R30 VGND.n0 VGND.t1 37.5
R31 VGND.n0 VGND.t0 36.818
R32 A1.n0 A1.t0 510.919
R33 A1.n0 A1.t1 200.832
R34 A1 A1.n0 93.69
R35 B1.n0 B1.t0 510.919
R36 B1.n0 B1.t1 199.226
R37 B1 B1.n0 51.974
C0 VPWR a_216_351# 0.04fF
C1 a_216_351# a_111_47# 0.02fF
C2 A1 VPWR 0.13fF
C3 A1 a_111_47# 0.10fF
C4 A2 a_216_351# 0.04fF
C5 A2 A1 0.08fF
C6 B1 VPWR 0.04fF
C7 B1 a_111_47# 0.01fF
C8 A2 B1 0.09fF
C9 A1 a_216_351# 0.00fF
C10 Y VPWR 0.38fF
C11 Y a_111_47# 0.05fF
C12 Y A2 0.03fF
C13 Y a_216_351# 0.02fF
C14 Y A1 0.00fF
C15 Y B1 0.21fF
C16 VPWR a_111_47# 0.01fF
C17 A2 VPWR 0.03fF
C18 A2 a_111_47# 0.11fF
.ends

