magic
tech sky130A
magscale 1 2
timestamp 1678746957
<< nwell >>
rect -38 315 866 998
<< nmos >>
rect 195 47 225 223
rect 349 47 379 223
rect 503 47 533 223
rect 657 47 687 223
<< pmos >>
rect 195 351 225 913
rect 349 351 379 913
rect 503 351 533 913
rect 657 351 687 913
<< ndiff >>
rect 115 173 195 223
rect 115 139 138 173
rect 172 139 195 173
rect 115 105 195 139
rect 115 71 138 105
rect 172 71 195 105
rect 115 47 195 71
rect 225 47 349 223
rect 379 173 503 223
rect 379 139 424 173
rect 458 139 503 173
rect 379 105 503 139
rect 379 71 424 105
rect 458 71 503 105
rect 379 47 503 71
rect 533 105 657 223
rect 533 71 544 105
rect 578 71 612 105
rect 646 71 657 105
rect 533 47 657 71
rect 687 173 767 223
rect 687 139 710 173
rect 744 139 767 173
rect 687 105 767 139
rect 687 71 710 105
rect 744 71 767 105
rect 687 47 767 71
<< pdiff >>
rect 115 889 195 913
rect 115 855 138 889
rect 172 855 195 889
rect 115 821 195 855
rect 115 787 138 821
rect 172 787 195 821
rect 115 753 195 787
rect 115 719 138 753
rect 172 719 195 753
rect 115 685 195 719
rect 115 651 138 685
rect 172 651 195 685
rect 115 617 195 651
rect 115 583 138 617
rect 172 583 195 617
rect 115 549 195 583
rect 115 515 138 549
rect 172 515 195 549
rect 115 481 195 515
rect 115 447 138 481
rect 172 447 195 481
rect 115 351 195 447
rect 225 889 349 913
rect 225 855 236 889
rect 270 855 304 889
rect 338 855 349 889
rect 225 821 349 855
rect 225 787 236 821
rect 270 787 304 821
rect 338 787 349 821
rect 225 753 349 787
rect 225 719 236 753
rect 270 719 304 753
rect 338 719 349 753
rect 225 685 349 719
rect 225 651 236 685
rect 270 651 304 685
rect 338 651 349 685
rect 225 617 349 651
rect 225 583 236 617
rect 270 583 304 617
rect 338 583 349 617
rect 225 549 349 583
rect 225 515 236 549
rect 270 515 304 549
rect 338 515 349 549
rect 225 351 349 515
rect 379 889 503 913
rect 379 855 424 889
rect 458 855 503 889
rect 379 821 503 855
rect 379 787 424 821
rect 458 787 503 821
rect 379 753 503 787
rect 379 719 424 753
rect 458 719 503 753
rect 379 685 503 719
rect 379 651 424 685
rect 458 651 503 685
rect 379 617 503 651
rect 379 583 424 617
rect 458 583 503 617
rect 379 549 503 583
rect 379 515 424 549
rect 458 515 503 549
rect 379 481 503 515
rect 379 447 424 481
rect 458 447 503 481
rect 379 351 503 447
rect 533 351 657 913
rect 687 891 767 913
rect 687 857 710 891
rect 744 857 767 891
rect 687 823 767 857
rect 687 789 710 823
rect 744 789 767 823
rect 687 755 767 789
rect 687 721 710 755
rect 744 721 767 755
rect 687 687 767 721
rect 687 653 710 687
rect 744 653 767 687
rect 687 619 767 653
rect 687 585 710 619
rect 744 585 767 619
rect 687 551 767 585
rect 687 517 710 551
rect 744 517 767 551
rect 687 483 767 517
rect 687 449 710 483
rect 744 449 767 483
rect 687 351 767 449
<< ndiffc >>
rect 138 139 172 173
rect 138 71 172 105
rect 424 139 458 173
rect 424 71 458 105
rect 544 71 578 105
rect 612 71 646 105
rect 710 139 744 173
rect 710 71 744 105
<< pdiffc >>
rect 138 855 172 889
rect 138 787 172 821
rect 138 719 172 753
rect 138 651 172 685
rect 138 583 172 617
rect 138 515 172 549
rect 138 447 172 481
rect 236 855 270 889
rect 304 855 338 889
rect 236 787 270 821
rect 304 787 338 821
rect 236 719 270 753
rect 304 719 338 753
rect 236 651 270 685
rect 304 651 338 685
rect 236 583 270 617
rect 304 583 338 617
rect 236 515 270 549
rect 304 515 338 549
rect 424 855 458 889
rect 424 787 458 821
rect 424 719 458 753
rect 424 651 458 685
rect 424 583 458 617
rect 424 515 458 549
rect 424 447 458 481
rect 710 857 744 891
rect 710 789 744 823
rect 710 721 744 755
rect 710 653 744 687
rect 710 585 744 619
rect 710 517 744 551
rect 710 449 744 483
<< psubdiff >>
rect 36 173 115 223
rect 36 139 58 173
rect 92 139 115 173
rect 36 105 115 139
rect 36 71 58 105
rect 92 71 115 105
rect 36 47 115 71
<< nsubdiff >>
rect 36 889 115 913
rect 36 855 59 889
rect 93 855 115 889
rect 36 821 115 855
rect 36 787 59 821
rect 93 787 115 821
rect 36 753 115 787
rect 36 719 59 753
rect 93 719 115 753
rect 36 685 115 719
rect 36 651 59 685
rect 93 651 115 685
rect 36 617 115 651
rect 36 583 59 617
rect 93 583 115 617
rect 36 549 115 583
rect 36 515 59 549
rect 93 515 115 549
rect 36 481 115 515
rect 36 447 59 481
rect 93 447 115 481
rect 36 351 115 447
<< psubdiffcont >>
rect 58 139 92 173
rect 58 71 92 105
<< nsubdiffcont >>
rect 59 855 93 889
rect 59 787 93 821
rect 59 719 93 753
rect 59 651 93 685
rect 59 583 93 617
rect 59 515 93 549
rect 59 447 93 481
<< poly >>
rect 195 913 225 939
rect 349 913 379 939
rect 503 913 533 939
rect 657 913 687 939
rect 195 314 225 351
rect 349 314 379 351
rect 503 314 533 351
rect 657 314 687 351
rect 61 304 225 314
rect 61 270 77 304
rect 111 270 145 304
rect 179 270 225 304
rect 61 260 225 270
rect 267 304 401 314
rect 267 270 283 304
rect 317 270 351 304
rect 385 270 401 304
rect 267 260 401 270
rect 443 304 579 314
rect 443 270 459 304
rect 493 270 527 304
rect 561 270 579 304
rect 443 260 579 270
rect 657 304 797 314
rect 657 270 679 304
rect 713 270 747 304
rect 781 270 797 304
rect 657 260 797 270
rect 195 223 225 260
rect 349 223 379 260
rect 503 223 533 260
rect 657 223 687 260
rect 195 21 225 47
rect 349 21 379 47
rect 503 21 533 47
rect 657 21 687 47
<< polycont >>
rect 77 270 111 304
rect 145 270 179 304
rect 283 270 317 304
rect 351 270 385 304
rect 459 270 493 304
rect 527 270 561 304
rect 679 270 713 304
rect 747 270 781 304
<< locali >>
rect 0 943 28 977
rect 62 943 121 977
rect 155 943 213 977
rect 247 943 305 977
rect 339 943 397 977
rect 431 943 489 977
rect 523 943 581 977
rect 615 943 673 977
rect 707 943 765 977
rect 799 943 828 977
rect 59 889 93 943
rect 59 821 93 855
rect 59 753 93 787
rect 59 685 93 719
rect 59 617 93 651
rect 59 549 93 583
rect 59 481 93 515
rect 59 431 93 447
rect 138 889 172 909
rect 138 821 172 855
rect 138 753 172 787
rect 138 685 172 719
rect 138 617 172 651
rect 138 549 172 583
rect 138 481 172 515
rect 236 889 339 943
rect 270 855 304 889
rect 338 855 339 889
rect 236 821 339 855
rect 270 787 304 821
rect 338 787 339 821
rect 236 753 339 787
rect 270 719 304 753
rect 338 719 339 753
rect 236 685 339 719
rect 270 651 304 685
rect 338 651 339 685
rect 236 617 339 651
rect 270 583 304 617
rect 338 583 339 617
rect 236 549 339 583
rect 270 515 304 549
rect 338 515 339 549
rect 236 499 339 515
rect 424 889 458 909
rect 424 821 458 855
rect 424 753 458 787
rect 424 685 458 719
rect 424 617 458 651
rect 424 549 458 583
rect 424 481 458 515
rect 172 447 424 465
rect 710 891 744 907
rect 710 823 744 857
rect 710 755 744 789
rect 744 721 745 730
rect 710 687 745 721
rect 744 653 745 687
rect 710 619 745 653
rect 744 585 745 619
rect 710 551 745 585
rect 744 517 745 551
rect 710 483 745 517
rect 138 431 458 447
rect 595 449 710 467
rect 744 449 745 483
rect 595 433 745 449
rect 77 304 179 383
rect 111 270 145 304
rect 77 254 179 270
rect 283 304 385 383
rect 317 270 351 304
rect 283 254 385 270
rect 459 304 561 383
rect 493 270 527 304
rect 459 254 561 270
rect 595 201 629 433
rect 678 304 781 383
rect 678 270 679 304
rect 713 270 747 304
rect 678 254 781 270
rect 58 173 184 190
rect 92 139 138 173
rect 172 139 184 173
rect 58 105 184 139
rect 92 71 138 105
rect 172 71 184 105
rect 58 17 184 71
rect 424 173 744 201
rect 458 166 710 173
rect 424 105 458 139
rect 710 105 744 139
rect 424 51 458 71
rect 527 71 544 105
rect 578 71 612 105
rect 646 71 662 105
rect 527 17 662 71
rect 710 51 744 71
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 28 943 62 977
rect 121 943 155 977
rect 213 943 247 977
rect 305 943 339 977
rect 397 943 431 977
rect 489 943 523 977
rect 581 943 615 977
rect 673 943 707 977
rect 765 943 799 977
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 977 828 1000
rect 0 943 28 977
rect 62 943 121 977
rect 155 943 213 977
rect 247 943 305 977
rect 339 943 397 977
rect 431 943 489 977
rect 523 943 581 977
rect 615 943 673 977
rect 707 943 765 977
rect 799 943 828 977
rect 0 920 828 943
rect 0 17 828 40
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -40 828 -17
<< labels >>
flabel locali s 121 343 155 377 0 FreeSans 240 0 0 0 A2
port 0 nsew signal input
flabel locali s 305 343 339 377 0 FreeSans 240 0 0 0 A1
port 1 nsew signal input
flabel locali s 489 343 523 377 0 FreeSans 240 0 0 0 B1
port 2 nsew signal input
flabel locali s 717 343 751 377 0 FreeSans 240 0 0 0 C1
port 3 nsew signal input
flabel metal1 s 397 943 431 977 0 FreeSans 240 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 397 -17 431 17 0 FreeSans 240 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 710 583 744 617 0 FreeSans 240 0 0 0 Y
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 960
string LEFclass CORE
string LEForigin 0 0
<< end >>
